
module progmem
(
// Closk & reset
input  wire         clk,
input  wire         rstn,

// PicoRV32 bus interface
input  wire         valid,
output wire         ready,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);

// ============================================================================

localparam  MEM_SIZE_BITS   = 12; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
localparam  MEM_ADDR_MASK   = 32'h0010_0000;

// ============================================================================

wire [MEM_SIZE_BITS-1:0]    mem_addr;
reg  [31:0]                 mem_data;

always @(posedge clk)
    case (mem_addr)

    'h0000: mem_data <= 32'h00000093;
    'h0001: mem_data <= 32'h00000193;
    'h0002: mem_data <= 32'h00000213;
    'h0003: mem_data <= 32'h00000293;
    'h0004: mem_data <= 32'h00000313;
    'h0005: mem_data <= 32'h00000393;
    'h0006: mem_data <= 32'h00000413;
    'h0007: mem_data <= 32'h00000493;
    'h0008: mem_data <= 32'h00000513;
    'h0009: mem_data <= 32'h00000593;
    'h000A: mem_data <= 32'h00000613;
    'h000B: mem_data <= 32'h00000693;
    'h000C: mem_data <= 32'h00000713;
    'h000D: mem_data <= 32'h00000793;
    'h000E: mem_data <= 32'h00000813;
    'h000F: mem_data <= 32'h00000893;
    'h0010: mem_data <= 32'h00000913;
    'h0011: mem_data <= 32'h00000993;
    'h0012: mem_data <= 32'h00000A13;
    'h0013: mem_data <= 32'h00000A93;
    'h0014: mem_data <= 32'h00000B13;
    'h0015: mem_data <= 32'h00000B93;
    'h0016: mem_data <= 32'h00000C13;
    'h0017: mem_data <= 32'h00000C93;
    'h0018: mem_data <= 32'h00000D13;
    'h0019: mem_data <= 32'h00000D93;
    'h001A: mem_data <= 32'h00000E13;
    'h001B: mem_data <= 32'h00000E93;
    'h001C: mem_data <= 32'h00000F13;
    'h001D: mem_data <= 32'h00000F93;
    'h001E: mem_data <= 32'h03000537;
    'h001F: mem_data <= 32'h00100593;
    'h0020: mem_data <= 32'h00B52023;
    'h0021: mem_data <= 32'h00000513;
    'h0022: mem_data <= 32'h00A52023;
    'h0023: mem_data <= 32'h00450513;
    'h0024: mem_data <= 32'hFE254CE3;
    'h0025: mem_data <= 32'h03000537;
    'h0026: mem_data <= 32'h00300593;
    'h0027: mem_data <= 32'h00B52023;
    'h0028: mem_data <= 32'h00003517;
    'h0029: mem_data <= 32'hC6C50513;
    'h002A: mem_data <= 32'h00000593;
    'h002B: mem_data <= 32'h00000613;
    'h002C: mem_data <= 32'h00C5DC63;
    'h002D: mem_data <= 32'h00052683;
    'h002E: mem_data <= 32'h00D5A023;
    'h002F: mem_data <= 32'h00450513;
    'h0030: mem_data <= 32'h00458593;
    'h0031: mem_data <= 32'hFEC5C8E3;
    'h0032: mem_data <= 32'h03000537;
    'h0033: mem_data <= 32'h00700593;
    'h0034: mem_data <= 32'h00B52023;
    'h0035: mem_data <= 32'h00000513;
    'h0036: mem_data <= 32'h00C00593;
    'h0037: mem_data <= 32'h00B55863;
    'h0038: mem_data <= 32'h00052023;
    'h0039: mem_data <= 32'h00450513;
    'h003A: mem_data <= 32'hFEB54CE3;
    'h003B: mem_data <= 32'h03000537;
    'h003C: mem_data <= 32'h00F00593;
    'h003D: mem_data <= 32'h00B52023;
    'h003E: mem_data <= 32'h045010EF;
    'h003F: mem_data <= 32'h0000006F;
    'h0040: mem_data <= 32'h020002B7;
    'h0041: mem_data <= 32'h12000313;
    'h0042: mem_data <= 32'h00629023;
    'h0043: mem_data <= 32'h000281A3;
    'h0044: mem_data <= 32'h02060863;
    'h0045: mem_data <= 32'h00800F13;
    'h0046: mem_data <= 32'h0FF67393;
    'h0047: mem_data <= 32'h0073DE93;
    'h0048: mem_data <= 32'h01D28023;
    'h0049: mem_data <= 32'h010EEE93;
    'h004A: mem_data <= 32'h01D28023;
    'h004B: mem_data <= 32'h00139393;
    'h004C: mem_data <= 32'h0FF3F393;
    'h004D: mem_data <= 32'hFFFF0F13;
    'h004E: mem_data <= 32'hFE0F12E3;
    'h004F: mem_data <= 32'h00628023;
    'h0050: mem_data <= 32'h04058663;
    'h0051: mem_data <= 32'h00800F13;
    'h0052: mem_data <= 32'h00054383;
    'h0053: mem_data <= 32'h0073DE93;
    'h0054: mem_data <= 32'h01D28023;
    'h0055: mem_data <= 32'h010EEE93;
    'h0056: mem_data <= 32'h01D28023;
    'h0057: mem_data <= 32'h0002CE83;
    'h0058: mem_data <= 32'h002EFE93;
    'h0059: mem_data <= 32'h001EDE93;
    'h005A: mem_data <= 32'h00139393;
    'h005B: mem_data <= 32'h01D3E3B3;
    'h005C: mem_data <= 32'h0FF3F393;
    'h005D: mem_data <= 32'hFFFF0F13;
    'h005E: mem_data <= 32'hFC0F1AE3;
    'h005F: mem_data <= 32'h00750023;
    'h0060: mem_data <= 32'h00150513;
    'h0061: mem_data <= 32'hFFF58593;
    'h0062: mem_data <= 32'hFB9FF06F;
    'h0063: mem_data <= 32'h08000313;
    'h0064: mem_data <= 32'h006281A3;
    'h0065: mem_data <= 32'h00008067;
    'h0066: mem_data <= 32'hFE010113;
    'h0067: mem_data <= 32'h00112E23;
    'h0068: mem_data <= 32'h00812C23;
    'h0069: mem_data <= 32'h02010413;
    'h006A: mem_data <= 32'h00050793;
    'h006B: mem_data <= 32'hFEF407A3;
    'h006C: mem_data <= 32'hFEF44703;
    'h006D: mem_data <= 32'h00A00793;
    'h006E: mem_data <= 32'h00F71663;
    'h006F: mem_data <= 32'h00D00513;
    'h0070: mem_data <= 32'hFD9FF0EF;
    'h0071: mem_data <= 32'h020007B7;
    'h0072: mem_data <= 32'h00878793;
    'h0073: mem_data <= 32'hFEF44703;
    'h0074: mem_data <= 32'h00E7A023;
    'h0075: mem_data <= 32'h00000013;
    'h0076: mem_data <= 32'h01C12083;
    'h0077: mem_data <= 32'h01812403;
    'h0078: mem_data <= 32'h02010113;
    'h0079: mem_data <= 32'h00008067;
    'h007A: mem_data <= 32'hFE010113;
    'h007B: mem_data <= 32'h00112E23;
    'h007C: mem_data <= 32'h00812C23;
    'h007D: mem_data <= 32'h02010413;
    'h007E: mem_data <= 32'hFEA42623;
    'h007F: mem_data <= 32'h01C0006F;
    'h0080: mem_data <= 32'hFEC42783;
    'h0081: mem_data <= 32'h00178713;
    'h0082: mem_data <= 32'hFEE42623;
    'h0083: mem_data <= 32'h0007C783;
    'h0084: mem_data <= 32'h00078513;
    'h0085: mem_data <= 32'hF85FF0EF;
    'h0086: mem_data <= 32'hFEC42783;
    'h0087: mem_data <= 32'h0007C783;
    'h0088: mem_data <= 32'hFE0790E3;
    'h0089: mem_data <= 32'h00000013;
    'h008A: mem_data <= 32'h00000013;
    'h008B: mem_data <= 32'h01C12083;
    'h008C: mem_data <= 32'h01812403;
    'h008D: mem_data <= 32'h02010113;
    'h008E: mem_data <= 32'h00008067;
    'h008F: mem_data <= 32'hFD010113;
    'h0090: mem_data <= 32'h02112623;
    'h0091: mem_data <= 32'h02812423;
    'h0092: mem_data <= 32'h03010413;
    'h0093: mem_data <= 32'hFCA42E23;
    'h0094: mem_data <= 32'hFCB42C23;
    'h0095: mem_data <= 32'h00700793;
    'h0096: mem_data <= 32'hFEF42623;
    'h0097: mem_data <= 32'h06C0006F;
    'h0098: mem_data <= 32'hFEC42783;
    'h0099: mem_data <= 32'h00279793;
    'h009A: mem_data <= 32'hFDC42703;
    'h009B: mem_data <= 32'h00F757B3;
    'h009C: mem_data <= 32'h00F7F793;
    'h009D: mem_data <= 32'h00102737;
    'h009E: mem_data <= 32'hA8470713;
    'h009F: mem_data <= 32'h00F707B3;
    'h00A0: mem_data <= 32'h0007C783;
    'h00A1: mem_data <= 32'hFEF405A3;
    'h00A2: mem_data <= 32'hFEB44703;
    'h00A3: mem_data <= 32'h03000793;
    'h00A4: mem_data <= 32'h00F71863;
    'h00A5: mem_data <= 32'hFEC42703;
    'h00A6: mem_data <= 32'hFD842783;
    'h00A7: mem_data <= 32'h00F75E63;
    'h00A8: mem_data <= 32'hFEB44783;
    'h00A9: mem_data <= 32'h00078513;
    'h00AA: mem_data <= 32'hEF1FF0EF;
    'h00AB: mem_data <= 32'hFEC42783;
    'h00AC: mem_data <= 32'hFCF42C23;
    'h00AD: mem_data <= 32'h0080006F;
    'h00AE: mem_data <= 32'h00000013;
    'h00AF: mem_data <= 32'hFEC42783;
    'h00B0: mem_data <= 32'hFFF78793;
    'h00B1: mem_data <= 32'hFEF42623;
    'h00B2: mem_data <= 32'hFEC42783;
    'h00B3: mem_data <= 32'hF807DAE3;
    'h00B4: mem_data <= 32'h00000013;
    'h00B5: mem_data <= 32'h00000013;
    'h00B6: mem_data <= 32'h02C12083;
    'h00B7: mem_data <= 32'h02812403;
    'h00B8: mem_data <= 32'h03010113;
    'h00B9: mem_data <= 32'h00008067;
    'h00BA: mem_data <= 32'hFE010113;
    'h00BB: mem_data <= 32'h00112E23;
    'h00BC: mem_data <= 32'h00812C23;
    'h00BD: mem_data <= 32'h02010413;
    'h00BE: mem_data <= 32'hFEA42623;
    'h00BF: mem_data <= 32'hFEC42703;
    'h00C0: mem_data <= 32'h06300793;
    'h00C1: mem_data <= 32'h00E7FA63;
    'h00C2: mem_data <= 32'h001027B7;
    'h00C3: mem_data <= 32'hA9878513;
    'h00C4: mem_data <= 32'hED9FF0EF;
    'h00C5: mem_data <= 32'h28C0006F;
    'h00C6: mem_data <= 32'hFEC42703;
    'h00C7: mem_data <= 32'h05900793;
    'h00C8: mem_data <= 32'h00E7FE63;
    'h00C9: mem_data <= 32'h03900513;
    'h00CA: mem_data <= 32'hE71FF0EF;
    'h00CB: mem_data <= 32'hFEC42783;
    'h00CC: mem_data <= 32'hFA678793;
    'h00CD: mem_data <= 32'hFEF42623;
    'h00CE: mem_data <= 32'h1200006F;
    'h00CF: mem_data <= 32'hFEC42703;
    'h00D0: mem_data <= 32'h04F00793;
    'h00D1: mem_data <= 32'h00E7FE63;
    'h00D2: mem_data <= 32'h03800513;
    'h00D3: mem_data <= 32'hE4DFF0EF;
    'h00D4: mem_data <= 32'hFEC42783;
    'h00D5: mem_data <= 32'hFB078793;
    'h00D6: mem_data <= 32'hFEF42623;
    'h00D7: mem_data <= 32'h0FC0006F;
    'h00D8: mem_data <= 32'hFEC42703;
    'h00D9: mem_data <= 32'h04500793;
    'h00DA: mem_data <= 32'h00E7FE63;
    'h00DB: mem_data <= 32'h03700513;
    'h00DC: mem_data <= 32'hE29FF0EF;
    'h00DD: mem_data <= 32'hFEC42783;
    'h00DE: mem_data <= 32'hFBA78793;
    'h00DF: mem_data <= 32'hFEF42623;
    'h00E0: mem_data <= 32'h0D80006F;
    'h00E1: mem_data <= 32'hFEC42703;
    'h00E2: mem_data <= 32'h03B00793;
    'h00E3: mem_data <= 32'h00E7FE63;
    'h00E4: mem_data <= 32'h03600513;
    'h00E5: mem_data <= 32'hE05FF0EF;
    'h00E6: mem_data <= 32'hFEC42783;
    'h00E7: mem_data <= 32'hFC478793;
    'h00E8: mem_data <= 32'hFEF42623;
    'h00E9: mem_data <= 32'h0B40006F;
    'h00EA: mem_data <= 32'hFEC42703;
    'h00EB: mem_data <= 32'h03100793;
    'h00EC: mem_data <= 32'h00E7FE63;
    'h00ED: mem_data <= 32'h03500513;
    'h00EE: mem_data <= 32'hDE1FF0EF;
    'h00EF: mem_data <= 32'hFEC42783;
    'h00F0: mem_data <= 32'hFCE78793;
    'h00F1: mem_data <= 32'hFEF42623;
    'h00F2: mem_data <= 32'h0900006F;
    'h00F3: mem_data <= 32'hFEC42703;
    'h00F4: mem_data <= 32'h02700793;
    'h00F5: mem_data <= 32'h00E7FE63;
    'h00F6: mem_data <= 32'h03400513;
    'h00F7: mem_data <= 32'hDBDFF0EF;
    'h00F8: mem_data <= 32'hFEC42783;
    'h00F9: mem_data <= 32'hFD878793;
    'h00FA: mem_data <= 32'hFEF42623;
    'h00FB: mem_data <= 32'h06C0006F;
    'h00FC: mem_data <= 32'hFEC42703;
    'h00FD: mem_data <= 32'h01D00793;
    'h00FE: mem_data <= 32'h00E7FE63;
    'h00FF: mem_data <= 32'h03300513;
    'h0100: mem_data <= 32'hD99FF0EF;
    'h0101: mem_data <= 32'hFEC42783;
    'h0102: mem_data <= 32'hFE278793;
    'h0103: mem_data <= 32'hFEF42623;
    'h0104: mem_data <= 32'h0480006F;
    'h0105: mem_data <= 32'hFEC42703;
    'h0106: mem_data <= 32'h01300793;
    'h0107: mem_data <= 32'h00E7FE63;
    'h0108: mem_data <= 32'h03200513;
    'h0109: mem_data <= 32'hD75FF0EF;
    'h010A: mem_data <= 32'hFEC42783;
    'h010B: mem_data <= 32'hFEC78793;
    'h010C: mem_data <= 32'hFEF42623;
    'h010D: mem_data <= 32'h0240006F;
    'h010E: mem_data <= 32'hFEC42703;
    'h010F: mem_data <= 32'h00900793;
    'h0110: mem_data <= 32'h00E7FC63;
    'h0111: mem_data <= 32'h03100513;
    'h0112: mem_data <= 32'hD51FF0EF;
    'h0113: mem_data <= 32'hFEC42783;
    'h0114: mem_data <= 32'hFF678793;
    'h0115: mem_data <= 32'hFEF42623;
    'h0116: mem_data <= 32'hFEC42703;
    'h0117: mem_data <= 32'h00800793;
    'h0118: mem_data <= 32'h00E7FE63;
    'h0119: mem_data <= 32'h03900513;
    'h011A: mem_data <= 32'hD31FF0EF;
    'h011B: mem_data <= 32'hFEC42783;
    'h011C: mem_data <= 32'hFF778793;
    'h011D: mem_data <= 32'hFEF42623;
    'h011E: mem_data <= 32'h1280006F;
    'h011F: mem_data <= 32'hFEC42703;
    'h0120: mem_data <= 32'h00700793;
    'h0121: mem_data <= 32'h00E7FE63;
    'h0122: mem_data <= 32'h03800513;
    'h0123: mem_data <= 32'hD0DFF0EF;
    'h0124: mem_data <= 32'hFEC42783;
    'h0125: mem_data <= 32'hFF878793;
    'h0126: mem_data <= 32'hFEF42623;
    'h0127: mem_data <= 32'h1040006F;
    'h0128: mem_data <= 32'hFEC42703;
    'h0129: mem_data <= 32'h00600793;
    'h012A: mem_data <= 32'h00E7FE63;
    'h012B: mem_data <= 32'h03700513;
    'h012C: mem_data <= 32'hCE9FF0EF;
    'h012D: mem_data <= 32'hFEC42783;
    'h012E: mem_data <= 32'hFF978793;
    'h012F: mem_data <= 32'hFEF42623;
    'h0130: mem_data <= 32'h0E00006F;
    'h0131: mem_data <= 32'hFEC42703;
    'h0132: mem_data <= 32'h00500793;
    'h0133: mem_data <= 32'h00E7FE63;
    'h0134: mem_data <= 32'h03600513;
    'h0135: mem_data <= 32'hCC5FF0EF;
    'h0136: mem_data <= 32'hFEC42783;
    'h0137: mem_data <= 32'hFFA78793;
    'h0138: mem_data <= 32'hFEF42623;
    'h0139: mem_data <= 32'h0BC0006F;
    'h013A: mem_data <= 32'hFEC42703;
    'h013B: mem_data <= 32'h00400793;
    'h013C: mem_data <= 32'h00E7FE63;
    'h013D: mem_data <= 32'h03500513;
    'h013E: mem_data <= 32'hCA1FF0EF;
    'h013F: mem_data <= 32'hFEC42783;
    'h0140: mem_data <= 32'hFFB78793;
    'h0141: mem_data <= 32'hFEF42623;
    'h0142: mem_data <= 32'h0980006F;
    'h0143: mem_data <= 32'hFEC42703;
    'h0144: mem_data <= 32'h00300793;
    'h0145: mem_data <= 32'h00E7FE63;
    'h0146: mem_data <= 32'h03400513;
    'h0147: mem_data <= 32'hC7DFF0EF;
    'h0148: mem_data <= 32'hFEC42783;
    'h0149: mem_data <= 32'hFFC78793;
    'h014A: mem_data <= 32'hFEF42623;
    'h014B: mem_data <= 32'h0740006F;
    'h014C: mem_data <= 32'hFEC42703;
    'h014D: mem_data <= 32'h00200793;
    'h014E: mem_data <= 32'h00E7FE63;
    'h014F: mem_data <= 32'h03300513;
    'h0150: mem_data <= 32'hC59FF0EF;
    'h0151: mem_data <= 32'hFEC42783;
    'h0152: mem_data <= 32'hFFD78793;
    'h0153: mem_data <= 32'hFEF42623;
    'h0154: mem_data <= 32'h0500006F;
    'h0155: mem_data <= 32'hFEC42703;
    'h0156: mem_data <= 32'h00100793;
    'h0157: mem_data <= 32'h00E7FE63;
    'h0158: mem_data <= 32'h03200513;
    'h0159: mem_data <= 32'hC35FF0EF;
    'h015A: mem_data <= 32'hFEC42783;
    'h015B: mem_data <= 32'hFFE78793;
    'h015C: mem_data <= 32'hFEF42623;
    'h015D: mem_data <= 32'h02C0006F;
    'h015E: mem_data <= 32'hFEC42783;
    'h015F: mem_data <= 32'h00078E63;
    'h0160: mem_data <= 32'h03100513;
    'h0161: mem_data <= 32'hC15FF0EF;
    'h0162: mem_data <= 32'hFEC42783;
    'h0163: mem_data <= 32'hFFF78793;
    'h0164: mem_data <= 32'hFEF42623;
    'h0165: mem_data <= 32'h00C0006F;
    'h0166: mem_data <= 32'h03000513;
    'h0167: mem_data <= 32'hBFDFF0EF;
    'h0168: mem_data <= 32'h01C12083;
    'h0169: mem_data <= 32'h01812403;
    'h016A: mem_data <= 32'h02010113;
    'h016B: mem_data <= 32'h00008067;
    'h016C: mem_data <= 32'hFD010113;
    'h016D: mem_data <= 32'h02112623;
    'h016E: mem_data <= 32'h02812423;
    'h016F: mem_data <= 32'h03010413;
    'h0170: mem_data <= 32'hFCA42E23;
    'h0171: mem_data <= 32'hFFF00793;
    'h0172: mem_data <= 32'hFEF42623;
    'h0173: mem_data <= 32'hC00027F3;
    'h0174: mem_data <= 32'hFEF42423;
    'h0175: mem_data <= 32'hFDC42783;
    'h0176: mem_data <= 32'h06078063;
    'h0177: mem_data <= 32'hFDC42503;
    'h0178: mem_data <= 32'hC09FF0EF;
    'h0179: mem_data <= 32'h0540006F;
    'h017A: mem_data <= 32'hC00027F3;
    'h017B: mem_data <= 32'hFEF42223;
    'h017C: mem_data <= 32'hFE442703;
    'h017D: mem_data <= 32'hFE842783;
    'h017E: mem_data <= 32'h40F707B3;
    'h017F: mem_data <= 32'hFEF42023;
    'h0180: mem_data <= 32'hFE042703;
    'h0181: mem_data <= 32'h01C9C7B7;
    'h0182: mem_data <= 32'h38078793;
    'h0183: mem_data <= 32'h00E7FE63;
    'h0184: mem_data <= 32'hFDC42783;
    'h0185: mem_data <= 32'h00078663;
    'h0186: mem_data <= 32'hFDC42503;
    'h0187: mem_data <= 32'hBCDFF0EF;
    'h0188: mem_data <= 32'hFE442783;
    'h0189: mem_data <= 32'hFEF42423;
    'h018A: mem_data <= 32'h020007B7;
    'h018B: mem_data <= 32'h00878793;
    'h018C: mem_data <= 32'h0007A783;
    'h018D: mem_data <= 32'hFEF42623;
    'h018E: mem_data <= 32'hFEC42703;
    'h018F: mem_data <= 32'hFFF00793;
    'h0190: mem_data <= 32'hFAF704E3;
    'h0191: mem_data <= 32'hFEC42783;
    'h0192: mem_data <= 32'h0FF7F793;
    'h0193: mem_data <= 32'h00078513;
    'h0194: mem_data <= 32'h02C12083;
    'h0195: mem_data <= 32'h02812403;
    'h0196: mem_data <= 32'h03010113;
    'h0197: mem_data <= 32'h00008067;
    'h0198: mem_data <= 32'hFF010113;
    'h0199: mem_data <= 32'h00112623;
    'h019A: mem_data <= 32'h00812423;
    'h019B: mem_data <= 32'h01010413;
    'h019C: mem_data <= 32'h00000513;
    'h019D: mem_data <= 32'hF3DFF0EF;
    'h019E: mem_data <= 32'h00050793;
    'h019F: mem_data <= 32'h00078513;
    'h01A0: mem_data <= 32'h00C12083;
    'h01A1: mem_data <= 32'h00812403;
    'h01A2: mem_data <= 32'h01010113;
    'h01A3: mem_data <= 32'h00008067;
    'h01A4: mem_data <= 32'hFD010113;
    'h01A5: mem_data <= 32'h02812623;
    'h01A6: mem_data <= 32'h03010413;
    'h01A7: mem_data <= 32'hFCA42E23;
    'h01A8: mem_data <= 32'hFE042423;
    'h01A9: mem_data <= 32'hFE042623;
    'h01AA: mem_data <= 32'hC00027F3;
    'h01AB: mem_data <= 32'hFEF42223;
    'h01AC: mem_data <= 32'hFE842703;
    'h01AD: mem_data <= 32'hFDC42783;
    'h01AE: mem_data <= 32'h02F75E63;
    'h01AF: mem_data <= 32'h01C0006F;
    'h01B0: mem_data <= 32'hC00027F3;
    'h01B1: mem_data <= 32'hFEF42023;
    'h01B2: mem_data <= 32'hFE042703;
    'h01B3: mem_data <= 32'hFE442783;
    'h01B4: mem_data <= 32'h40F707B3;
    'h01B5: mem_data <= 32'hFEF42623;
    'h01B6: mem_data <= 32'hFEC42703;
    'h01B7: mem_data <= 32'h01C9C7B7;
    'h01B8: mem_data <= 32'h37F78793;
    'h01B9: mem_data <= 32'hFCE7FEE3;
    'h01BA: mem_data <= 32'hFE842783;
    'h01BB: mem_data <= 32'h00178793;
    'h01BC: mem_data <= 32'hFEF42423;
    'h01BD: mem_data <= 32'h00000013;
    'h01BE: mem_data <= 32'h02C12403;
    'h01BF: mem_data <= 32'h03010113;
    'h01C0: mem_data <= 32'h00008067;
    'h01C1: mem_data <= 32'hFE010113;
    'h01C2: mem_data <= 32'h00112E23;
    'h01C3: mem_data <= 32'h00812C23;
    'h01C4: mem_data <= 32'h02010413;
    'h01C5: mem_data <= 32'h030007B7;
    'h01C6: mem_data <= 32'h0007A023;
    'h01C7: mem_data <= 32'h06400793;
    'h01C8: mem_data <= 32'hFEF42623;
    'h01C9: mem_data <= 32'h1580006F;
    'h01CA: mem_data <= 32'h001027B7;
    'h01CB: mem_data <= 32'hAA078513;
    'h01CC: mem_data <= 32'hAB9FF0EF;
    'h01CD: mem_data <= 32'hF2DFF0EF;
    'h01CE: mem_data <= 32'h00050793;
    'h01CF: mem_data <= 32'hFEF405A3;
    'h01D0: mem_data <= 32'hFEB44703;
    'h01D1: mem_data <= 32'h02000793;
    'h01D2: mem_data <= 32'h00E7FE63;
    'h01D3: mem_data <= 32'hFEB44703;
    'h01D4: mem_data <= 32'h07E00793;
    'h01D5: mem_data <= 32'h00E7E863;
    'h01D6: mem_data <= 32'hFEB44783;
    'h01D7: mem_data <= 32'h00078513;
    'h01D8: mem_data <= 32'hA39FF0EF;
    'h01D9: mem_data <= 32'h001027B7;
    'h01DA: mem_data <= 32'hAD878513;
    'h01DB: mem_data <= 32'hA7DFF0EF;
    'h01DC: mem_data <= 32'hFEB44783;
    'h01DD: mem_data <= 32'hFCF78793;
    'h01DE: mem_data <= 32'h04100713;
    'h01DF: mem_data <= 32'h0EF76863;
    'h01E0: mem_data <= 32'h00279713;
    'h01E1: mem_data <= 32'h001027B7;
    'h01E2: mem_data <= 32'hADC78793;
    'h01E3: mem_data <= 32'h00F707B3;
    'h01E4: mem_data <= 32'h0007A783;
    'h01E5: mem_data <= 32'h00078067;
    'h01E6: mem_data <= 32'h030007B7;
    'h01E7: mem_data <= 32'h0007A703;
    'h01E8: mem_data <= 32'h030007B7;
    'h01E9: mem_data <= 32'h00174713;
    'h01EA: mem_data <= 32'h00E7A023;
    'h01EB: mem_data <= 32'h0C40006F;
    'h01EC: mem_data <= 32'h030007B7;
    'h01ED: mem_data <= 32'h0007A703;
    'h01EE: mem_data <= 32'h030007B7;
    'h01EF: mem_data <= 32'h00274713;
    'h01F0: mem_data <= 32'h00E7A023;
    'h01F1: mem_data <= 32'h0AC0006F;
    'h01F2: mem_data <= 32'h030007B7;
    'h01F3: mem_data <= 32'h0007A703;
    'h01F4: mem_data <= 32'h030007B7;
    'h01F5: mem_data <= 32'h00474713;
    'h01F6: mem_data <= 32'h00E7A023;
    'h01F7: mem_data <= 32'h0940006F;
    'h01F8: mem_data <= 32'h030007B7;
    'h01F9: mem_data <= 32'h0007A703;
    'h01FA: mem_data <= 32'h030007B7;
    'h01FB: mem_data <= 32'h00874713;
    'h01FC: mem_data <= 32'h00E7A023;
    'h01FD: mem_data <= 32'h07C0006F;
    'h01FE: mem_data <= 32'h030007B7;
    'h01FF: mem_data <= 32'h0007A703;
    'h0200: mem_data <= 32'h030007B7;
    'h0201: mem_data <= 32'h01074713;
    'h0202: mem_data <= 32'h00E7A023;
    'h0203: mem_data <= 32'h0640006F;
    'h0204: mem_data <= 32'h030007B7;
    'h0205: mem_data <= 32'h0007A703;
    'h0206: mem_data <= 32'h030007B7;
    'h0207: mem_data <= 32'h02074713;
    'h0208: mem_data <= 32'h00E7A023;
    'h0209: mem_data <= 32'h04C0006F;
    'h020A: mem_data <= 32'h030007B7;
    'h020B: mem_data <= 32'h0007A703;
    'h020C: mem_data <= 32'h030007B7;
    'h020D: mem_data <= 32'h04074713;
    'h020E: mem_data <= 32'h00E7A023;
    'h020F: mem_data <= 32'h0340006F;
    'h0210: mem_data <= 32'h030007B7;
    'h0211: mem_data <= 32'h0007A703;
    'h0212: mem_data <= 32'h030007B7;
    'h0213: mem_data <= 32'h08074713;
    'h0214: mem_data <= 32'h00E7A023;
    'h0215: mem_data <= 32'h01C0006F;
    'h0216: mem_data <= 32'h030007B7;
    'h0217: mem_data <= 32'h0007A023;
    'h0218: mem_data <= 32'h00000013;
    'h0219: mem_data <= 32'h21D000EF;
    'h021A: mem_data <= 32'h0200006F;
    'h021B: mem_data <= 32'h00000013;
    'h021C: mem_data <= 32'hFEC42783;
    'h021D: mem_data <= 32'hFFF78793;
    'h021E: mem_data <= 32'hFEF42623;
    'h021F: mem_data <= 32'hFEC42783;
    'h0220: mem_data <= 32'hEAF044E3;
    'h0221: mem_data <= 32'h00000013;
    'h0222: mem_data <= 32'h00000013;
    'h0223: mem_data <= 32'h01C12083;
    'h0224: mem_data <= 32'h01812403;
    'h0225: mem_data <= 32'h02010113;
    'h0226: mem_data <= 32'h00008067;
    'h0227: mem_data <= 32'hFF010113;
    'h0228: mem_data <= 32'h00112623;
    'h0229: mem_data <= 32'h00812423;
    'h022A: mem_data <= 32'h01010413;
    'h022B: mem_data <= 32'h001027B7;
    'h022C: mem_data <= 32'hBE478513;
    'h022D: mem_data <= 32'h935FF0EF;
    'h022E: mem_data <= 32'h030007B7;
    'h022F: mem_data <= 32'h10078793;
    'h0230: mem_data <= 32'h0007A783;
    'h0231: mem_data <= 32'h1007F713;
    'h0232: mem_data <= 32'h10000793;
    'h0233: mem_data <= 32'h00F71A63;
    'h0234: mem_data <= 32'h001027B7;
    'h0235: mem_data <= 32'hBF078513;
    'h0236: mem_data <= 32'h911FF0EF;
    'h0237: mem_data <= 32'h0100006F;
    'h0238: mem_data <= 32'h001027B7;
    'h0239: mem_data <= 32'hBF878513;
    'h023A: mem_data <= 32'h901FF0EF;
    'h023B: mem_data <= 32'h001027B7;
    'h023C: mem_data <= 32'hBFC78513;
    'h023D: mem_data <= 32'h8F5FF0EF;
    'h023E: mem_data <= 32'h030007B7;
    'h023F: mem_data <= 32'h10078793;
    'h0240: mem_data <= 32'h0007A783;
    'h0241: mem_data <= 32'h2007F713;
    'h0242: mem_data <= 32'h20000793;
    'h0243: mem_data <= 32'h00F71A63;
    'h0244: mem_data <= 32'h001027B7;
    'h0245: mem_data <= 32'hC0878513;
    'h0246: mem_data <= 32'h8D1FF0EF;
    'h0247: mem_data <= 32'h0100006F;
    'h0248: mem_data <= 32'h001027B7;
    'h0249: mem_data <= 32'hC1078513;
    'h024A: mem_data <= 32'h8C1FF0EF;
    'h024B: mem_data <= 32'h001027B7;
    'h024C: mem_data <= 32'hC1878513;
    'h024D: mem_data <= 32'h8B5FF0EF;
    'h024E: mem_data <= 32'h030007B7;
    'h024F: mem_data <= 32'h10078793;
    'h0250: mem_data <= 32'h0007A783;
    'h0251: mem_data <= 32'h0017F713;
    'h0252: mem_data <= 32'h00100793;
    'h0253: mem_data <= 32'h00F71A63;
    'h0254: mem_data <= 32'h001027B7;
    'h0255: mem_data <= 32'hBF078513;
    'h0256: mem_data <= 32'h891FF0EF;
    'h0257: mem_data <= 32'h0100006F;
    'h0258: mem_data <= 32'h001027B7;
    'h0259: mem_data <= 32'hBF878513;
    'h025A: mem_data <= 32'h881FF0EF;
    'h025B: mem_data <= 32'h001027B7;
    'h025C: mem_data <= 32'hC1878513;
    'h025D: mem_data <= 32'h875FF0EF;
    'h025E: mem_data <= 32'h030007B7;
    'h025F: mem_data <= 32'h10078793;
    'h0260: mem_data <= 32'h0007A783;
    'h0261: mem_data <= 32'h0027F713;
    'h0262: mem_data <= 32'h00200793;
    'h0263: mem_data <= 32'h00F71A63;
    'h0264: mem_data <= 32'h001027B7;
    'h0265: mem_data <= 32'hBF078513;
    'h0266: mem_data <= 32'h851FF0EF;
    'h0267: mem_data <= 32'h0100006F;
    'h0268: mem_data <= 32'h001027B7;
    'h0269: mem_data <= 32'hBF878513;
    'h026A: mem_data <= 32'h841FF0EF;
    'h026B: mem_data <= 32'h001027B7;
    'h026C: mem_data <= 32'hC1878513;
    'h026D: mem_data <= 32'h835FF0EF;
    'h026E: mem_data <= 32'h030007B7;
    'h026F: mem_data <= 32'h10078793;
    'h0270: mem_data <= 32'h0007A783;
    'h0271: mem_data <= 32'h0047F713;
    'h0272: mem_data <= 32'h00400793;
    'h0273: mem_data <= 32'h00F71A63;
    'h0274: mem_data <= 32'h001027B7;
    'h0275: mem_data <= 32'hBF078513;
    'h0276: mem_data <= 32'h811FF0EF;
    'h0277: mem_data <= 32'h0100006F;
    'h0278: mem_data <= 32'h001027B7;
    'h0279: mem_data <= 32'hBF878513;
    'h027A: mem_data <= 32'h801FF0EF;
    'h027B: mem_data <= 32'h001027B7;
    'h027C: mem_data <= 32'hC1878513;
    'h027D: mem_data <= 32'hFF4FF0EF;
    'h027E: mem_data <= 32'h030007B7;
    'h027F: mem_data <= 32'h10078793;
    'h0280: mem_data <= 32'h0007A783;
    'h0281: mem_data <= 32'h0087F713;
    'h0282: mem_data <= 32'h00800793;
    'h0283: mem_data <= 32'h00F71A63;
    'h0284: mem_data <= 32'h001027B7;
    'h0285: mem_data <= 32'hC0878513;
    'h0286: mem_data <= 32'hFD0FF0EF;
    'h0287: mem_data <= 32'h0100006F;
    'h0288: mem_data <= 32'h001027B7;
    'h0289: mem_data <= 32'hC1078513;
    'h028A: mem_data <= 32'hFC0FF0EF;
    'h028B: mem_data <= 32'h00000013;
    'h028C: mem_data <= 32'h00C12083;
    'h028D: mem_data <= 32'h00812403;
    'h028E: mem_data <= 32'h01010113;
    'h028F: mem_data <= 32'h00008067;
    'h0290: mem_data <= 32'hFF010113;
    'h0291: mem_data <= 32'h00812623;
    'h0292: mem_data <= 32'h01010413;
    'h0293: mem_data <= 32'h060107B7;
    'h0294: mem_data <= 32'h10078793;
    'h0295: mem_data <= 32'h0007A783;
    'h0296: mem_data <= 32'h0FF7F713;
    'h0297: mem_data <= 32'h00E00023;
    'h0298: mem_data <= 32'h0180006F;
    'h0299: mem_data <= 32'h060107B7;
    'h029A: mem_data <= 32'h10078793;
    'h029B: mem_data <= 32'h0007A783;
    'h029C: mem_data <= 32'h0FF7F713;
    'h029D: mem_data <= 32'h00E00023;
    'h029E: mem_data <= 32'h00004783;
    'h029F: mem_data <= 32'h0027F793;
    'h02A0: mem_data <= 32'hFE0792E3;
    'h02A1: mem_data <= 32'h00000013;
    'h02A2: mem_data <= 32'h00000013;
    'h02A3: mem_data <= 32'h00C12403;
    'h02A4: mem_data <= 32'h01010113;
    'h02A5: mem_data <= 32'h00008067;
    'h02A6: mem_data <= 32'hFE010113;
    'h02A7: mem_data <= 32'h00112E23;
    'h02A8: mem_data <= 32'h00812C23;
    'h02A9: mem_data <= 32'h02010413;
    'h02AA: mem_data <= 32'h00050793;
    'h02AB: mem_data <= 32'hFEF407A3;
    'h02AC: mem_data <= 32'h060007B7;
    'h02AD: mem_data <= 32'h30078793;
    'h02AE: mem_data <= 32'hFEF44703;
    'h02AF: mem_data <= 32'h00E7A023;
    'h02B0: mem_data <= 32'h060007B7;
    'h02B1: mem_data <= 32'h40078793;
    'h02B2: mem_data <= 32'h01000713;
    'h02B3: mem_data <= 32'h00E7A023;
    'h02B4: mem_data <= 32'hF71FF0EF;
    'h02B5: mem_data <= 32'h00000013;
    'h02B6: mem_data <= 32'h01C12083;
    'h02B7: mem_data <= 32'h01812403;
    'h02B8: mem_data <= 32'h02010113;
    'h02B9: mem_data <= 32'h00008067;
    'h02BA: mem_data <= 32'hFE010113;
    'h02BB: mem_data <= 32'h00112E23;
    'h02BC: mem_data <= 32'h00812C23;
    'h02BD: mem_data <= 32'h02010413;
    'h02BE: mem_data <= 32'h00050793;
    'h02BF: mem_data <= 32'h00058713;
    'h02C0: mem_data <= 32'hFEF407A3;
    'h02C1: mem_data <= 32'h00070793;
    'h02C2: mem_data <= 32'hFEF40723;
    'h02C3: mem_data <= 32'hFEE44783;
    'h02C4: mem_data <= 32'h00078E63;
    'h02C5: mem_data <= 32'hFEF44783;
    'h02C6: mem_data <= 32'h00179713;
    'h02C7: mem_data <= 32'h060007B7;
    'h02C8: mem_data <= 32'h30078793;
    'h02C9: mem_data <= 32'h00E7A023;
    'h02CA: mem_data <= 32'h01C0006F;
    'h02CB: mem_data <= 32'hFEF44783;
    'h02CC: mem_data <= 32'h00179793;
    'h02CD: mem_data <= 32'h0017E713;
    'h02CE: mem_data <= 32'h060007B7;
    'h02CF: mem_data <= 32'h30078793;
    'h02D0: mem_data <= 32'h00E7A023;
    'h02D1: mem_data <= 32'h060007B7;
    'h02D2: mem_data <= 32'h40078793;
    'h02D3: mem_data <= 32'h09000713;
    'h02D4: mem_data <= 32'h00E7A023;
    'h02D5: mem_data <= 32'hEEDFF0EF;
    'h02D6: mem_data <= 32'h00000013;
    'h02D7: mem_data <= 32'h01C12083;
    'h02D8: mem_data <= 32'h01812403;
    'h02D9: mem_data <= 32'h02010113;
    'h02DA: mem_data <= 32'h00008067;
    'h02DB: mem_data <= 32'hFF010113;
    'h02DC: mem_data <= 32'h00112623;
    'h02DD: mem_data <= 32'h00812423;
    'h02DE: mem_data <= 32'h01010413;
    'h02DF: mem_data <= 32'h060007B7;
    'h02E0: mem_data <= 32'h40078793;
    'h02E1: mem_data <= 32'h02000713;
    'h02E2: mem_data <= 32'h00E7A023;
    'h02E3: mem_data <= 32'hEB5FF0EF;
    'h02E4: mem_data <= 32'h00000013;
    'h02E5: mem_data <= 32'h00C12083;
    'h02E6: mem_data <= 32'h00812403;
    'h02E7: mem_data <= 32'h01010113;
    'h02E8: mem_data <= 32'h00008067;
    'h02E9: mem_data <= 32'hFF010113;
    'h02EA: mem_data <= 32'h00112623;
    'h02EB: mem_data <= 32'h00812423;
    'h02EC: mem_data <= 32'h01010413;
    'h02ED: mem_data <= 32'h060007B7;
    'h02EE: mem_data <= 32'h40078793;
    'h02EF: mem_data <= 32'h04800713;
    'h02F0: mem_data <= 32'h00E7A023;
    'h02F1: mem_data <= 32'hE7DFF0EF;
    'h02F2: mem_data <= 32'h00000013;
    'h02F3: mem_data <= 32'h00C12083;
    'h02F4: mem_data <= 32'h00812403;
    'h02F5: mem_data <= 32'h01010113;
    'h02F6: mem_data <= 32'h00008067;
    'h02F7: mem_data <= 32'hFD010113;
    'h02F8: mem_data <= 32'h02112623;
    'h02F9: mem_data <= 32'h02812423;
    'h02FA: mem_data <= 32'h03010413;
    'h02FB: mem_data <= 32'h00050793;
    'h02FC: mem_data <= 32'hFCF40FA3;
    'h02FD: mem_data <= 32'hFE0407A3;
    'h02FE: mem_data <= 32'hDDCCC7B7;
    'h02FF: mem_data <= 32'hBAA78793;
    'h0300: mem_data <= 32'hFEF42423;
    'h0301: mem_data <= 32'h001027B7;
    'h0302: mem_data <= 32'hC2478513;
    'h0303: mem_data <= 32'hDDCFF0EF;
    'h0304: mem_data <= 32'h001027B7;
    'h0305: mem_data <= 32'hC3C78513;
    'h0306: mem_data <= 32'hDD0FF0EF;
    'h0307: mem_data <= 32'h001027B7;
    'h0308: mem_data <= 32'hC4878513;
    'h0309: mem_data <= 32'hDC4FF0EF;
    'h030A: mem_data <= 32'h060007B7;
    'h030B: mem_data <= 32'hFDF44703;
    'h030C: mem_data <= 32'h00E7A023;
    'h030D: mem_data <= 32'h060007B7;
    'h030E: mem_data <= 32'h10078793;
    'h030F: mem_data <= 32'h0007A023;
    'h0310: mem_data <= 32'h060007B7;
    'h0311: mem_data <= 32'h20078793;
    'h0312: mem_data <= 32'h08000713;
    'h0313: mem_data <= 32'h00E7A023;
    'h0314: mem_data <= 32'h00100593;
    'h0315: mem_data <= 32'h01000513;
    'h0316: mem_data <= 32'hE91FF0EF;
    'h0317: mem_data <= 32'h00000513;
    'h0318: mem_data <= 32'hE39FF0EF;
    'h0319: mem_data <= 32'h001027B7;
    'h031A: mem_data <= 32'hC6078513;
    'h031B: mem_data <= 32'hD7CFF0EF;
    'h031C: mem_data <= 32'h00A00513;
    'h031D: mem_data <= 32'hA1DFF0EF;
    'h031E: mem_data <= 32'h000002A3;
    'h031F: mem_data <= 32'h05C0006F;
    'h0320: mem_data <= 32'h00504783;
    'h0321: mem_data <= 32'hFF078793;
    'h0322: mem_data <= 32'h008787B3;
    'h0323: mem_data <= 32'hFF87C783;
    'h0324: mem_data <= 32'h00078513;
    'h0325: mem_data <= 32'hE05FF0EF;
    'h0326: mem_data <= 32'h00504783;
    'h0327: mem_data <= 32'hFF078793;
    'h0328: mem_data <= 32'h008787B3;
    'h0329: mem_data <= 32'hFF87C783;
    'h032A: mem_data <= 32'h00200593;
    'h032B: mem_data <= 32'h00078513;
    'h032C: mem_data <= 32'hD8CFF0EF;
    'h032D: mem_data <= 32'h001027B7;
    'h032E: mem_data <= 32'hC6C78513;
    'h032F: mem_data <= 32'hD2CFF0EF;
    'h0330: mem_data <= 32'h00A00513;
    'h0331: mem_data <= 32'h9CDFF0EF;
    'h0332: mem_data <= 32'h00504783;
    'h0333: mem_data <= 32'h00178793;
    'h0334: mem_data <= 32'h0FF7F713;
    'h0335: mem_data <= 32'h00E002A3;
    'h0336: mem_data <= 32'h00504703;
    'h0337: mem_data <= 32'h00300793;
    'h0338: mem_data <= 32'hFAE7F0E3;
    'h0339: mem_data <= 32'hEC1FF0EF;
    'h033A: mem_data <= 32'h00A00513;
    'h033B: mem_data <= 32'h9A5FF0EF;
    'h033C: mem_data <= 32'h001027B7;
    'h033D: mem_data <= 32'hC7078513;
    'h033E: mem_data <= 32'hCF0FF0EF;
    'h033F: mem_data <= 32'h00A00513;
    'h0340: mem_data <= 32'h991FF0EF;
    'h0341: mem_data <= 32'h000002A3;
    'h0342: mem_data <= 32'h0940006F;
    'h0343: mem_data <= 32'h00100593;
    'h0344: mem_data <= 32'h01000513;
    'h0345: mem_data <= 32'hDD5FF0EF;
    'h0346: mem_data <= 32'h00504783;
    'h0347: mem_data <= 32'h00078513;
    'h0348: mem_data <= 32'hD79FF0EF;
    'h0349: mem_data <= 32'h00000593;
    'h034A: mem_data <= 32'h01000513;
    'h034B: mem_data <= 32'hDBDFF0EF;
    'h034C: mem_data <= 32'hE3DFF0EF;
    'h034D: mem_data <= 32'h060107B7;
    'h034E: mem_data <= 32'h0007A783;
    'h034F: mem_data <= 32'hFEF40723;
    'h0350: mem_data <= 32'h00504783;
    'h0351: mem_data <= 32'hFF078793;
    'h0352: mem_data <= 32'h008787B3;
    'h0353: mem_data <= 32'hFF87C783;
    'h0354: mem_data <= 32'hFEE44703;
    'h0355: mem_data <= 32'h00F71863;
    'h0356: mem_data <= 32'hFEF44783;
    'h0357: mem_data <= 32'h00178793;
    'h0358: mem_data <= 32'hFEF407A3;
    'h0359: mem_data <= 32'hFEE44783;
    'h035A: mem_data <= 32'h00200593;
    'h035B: mem_data <= 32'h00078513;
    'h035C: mem_data <= 32'hCCCFF0EF;
    'h035D: mem_data <= 32'h001027B7;
    'h035E: mem_data <= 32'hC6C78513;
    'h035F: mem_data <= 32'hC6CFF0EF;
    'h0360: mem_data <= 32'hE25FF0EF;
    'h0361: mem_data <= 32'h00A00513;
    'h0362: mem_data <= 32'h909FF0EF;
    'h0363: mem_data <= 32'h00504783;
    'h0364: mem_data <= 32'h00178793;
    'h0365: mem_data <= 32'h0FF7F713;
    'h0366: mem_data <= 32'h00E002A3;
    'h0367: mem_data <= 32'h00504703;
    'h0368: mem_data <= 32'h00300793;
    'h0369: mem_data <= 32'hF6E7F4E3;
    'h036A: mem_data <= 32'hFEF44703;
    'h036B: mem_data <= 32'h00400793;
    'h036C: mem_data <= 32'h00F71A63;
    'h036D: mem_data <= 32'h001027B7;
    'h036E: mem_data <= 32'hC7C78513;
    'h036F: mem_data <= 32'hC2CFF0EF;
    'h0370: mem_data <= 32'h0100006F;
    'h0371: mem_data <= 32'h001027B7;
    'h0372: mem_data <= 32'hC9078513;
    'h0373: mem_data <= 32'hC1CFF0EF;
    'h0374: mem_data <= 32'h00000013;
    'h0375: mem_data <= 32'h02C12083;
    'h0376: mem_data <= 32'h02812403;
    'h0377: mem_data <= 32'h03010113;
    'h0378: mem_data <= 32'h00008067;
    'h0379: mem_data <= 32'hFF010113;
    'h037A: mem_data <= 32'h00812623;
    'h037B: mem_data <= 32'h01010413;
    'h037C: mem_data <= 32'h050107B7;
    'h037D: mem_data <= 32'h10078793;
    'h037E: mem_data <= 32'h0007A783;
    'h037F: mem_data <= 32'h0FF7F713;
    'h0380: mem_data <= 32'h00E000A3;
    'h0381: mem_data <= 32'h02C0006F;
    'h0382: mem_data <= 32'h050107B7;
    'h0383: mem_data <= 32'h10078793;
    'h0384: mem_data <= 32'h0007A783;
    'h0385: mem_data <= 32'h0FF7F713;
    'h0386: mem_data <= 32'h00E000A3;
    'h0387: mem_data <= 32'h050107B7;
    'h0388: mem_data <= 32'h10078793;
    'h0389: mem_data <= 32'h0007A783;
    'h038A: mem_data <= 32'h0FF7F713;
    'h038B: mem_data <= 32'h00E000A3;
    'h038C: mem_data <= 32'h00104783;
    'h038D: mem_data <= 32'h0027F793;
    'h038E: mem_data <= 32'hFC0798E3;
    'h038F: mem_data <= 32'h00000013;
    'h0390: mem_data <= 32'h00000013;
    'h0391: mem_data <= 32'h00C12403;
    'h0392: mem_data <= 32'h01010113;
    'h0393: mem_data <= 32'h00008067;
    'h0394: mem_data <= 32'hFF010113;
    'h0395: mem_data <= 32'h00812623;
    'h0396: mem_data <= 32'h01010413;
    'h0397: mem_data <= 32'h050107B7;
    'h0398: mem_data <= 32'h10078793;
    'h0399: mem_data <= 32'h0007A783;
    'h039A: mem_data <= 32'h0FF7F713;
    'h039B: mem_data <= 32'h00E000A3;
    'h039C: mem_data <= 32'h02C0006F;
    'h039D: mem_data <= 32'h050107B7;
    'h039E: mem_data <= 32'h10078793;
    'h039F: mem_data <= 32'h0007A783;
    'h03A0: mem_data <= 32'h0FF7F713;
    'h03A1: mem_data <= 32'h00E000A3;
    'h03A2: mem_data <= 32'h050107B7;
    'h03A3: mem_data <= 32'h10078793;
    'h03A4: mem_data <= 32'h0007A783;
    'h03A5: mem_data <= 32'h0FF7F713;
    'h03A6: mem_data <= 32'h00E000A3;
    'h03A7: mem_data <= 32'h00104783;
    'h03A8: mem_data <= 32'h0017F793;
    'h03A9: mem_data <= 32'hFC0788E3;
    'h03AA: mem_data <= 32'h00000013;
    'h03AB: mem_data <= 32'h00000013;
    'h03AC: mem_data <= 32'h00C12403;
    'h03AD: mem_data <= 32'h01010113;
    'h03AE: mem_data <= 32'h00008067;
    'h03AF: mem_data <= 32'hFE010113;
    'h03B0: mem_data <= 32'h00112E23;
    'h03B1: mem_data <= 32'h00812C23;
    'h03B2: mem_data <= 32'h02010413;
    'h03B3: mem_data <= 32'h00050793;
    'h03B4: mem_data <= 32'hFEF407A3;
    'h03B5: mem_data <= 32'h050007B7;
    'h03B6: mem_data <= 32'h20078793;
    'h03B7: mem_data <= 32'hFEF44703;
    'h03B8: mem_data <= 32'h00E7A023;
    'h03B9: mem_data <= 32'hF01FF0EF;
    'h03BA: mem_data <= 32'h00000013;
    'h03BB: mem_data <= 32'h01C12083;
    'h03BC: mem_data <= 32'h01812403;
    'h03BD: mem_data <= 32'h02010113;
    'h03BE: mem_data <= 32'h00008067;
    'h03BF: mem_data <= 32'hFC010113;
    'h03C0: mem_data <= 32'h02112E23;
    'h03C1: mem_data <= 32'h02812C23;
    'h03C2: mem_data <= 32'h04010413;
    'h03C3: mem_data <= 32'h00050793;
    'h03C4: mem_data <= 32'hFCF407A3;
    'h03C5: mem_data <= 32'hFE0407A3;
    'h03C6: mem_data <= 32'h001027B7;
    'h03C7: mem_data <= 32'hC2478513;
    'h03C8: mem_data <= 32'hAC8FF0EF;
    'h03C9: mem_data <= 32'h001027B7;
    'h03CA: mem_data <= 32'hCA878513;
    'h03CB: mem_data <= 32'hABCFF0EF;
    'h03CC: mem_data <= 32'h001027B7;
    'h03CD: mem_data <= 32'hC4878513;
    'h03CE: mem_data <= 32'hAB0FF0EF;
    'h03CF: mem_data <= 32'h050007B7;
    'h03D0: mem_data <= 32'h30078793;
    'h03D1: mem_data <= 32'h0007A023;
    'h03D2: mem_data <= 32'h00000123;
    'h03D3: mem_data <= 32'h2D00006F;
    'h03D4: mem_data <= 32'h000001A3;
    'h03D5: mem_data <= 32'h2AC0006F;
    'h03D6: mem_data <= 32'h050007B7;
    'h03D7: mem_data <= 32'h30078793;
    'h03D8: mem_data <= 32'h00100713;
    'h03D9: mem_data <= 32'h00E7A023;
    'h03DA: mem_data <= 32'h001027B7;
    'h03DB: mem_data <= 32'hCB478513;
    'h03DC: mem_data <= 32'hA78FF0EF;
    'h03DD: mem_data <= 32'h00204783;
    'h03DE: mem_data <= 32'h00078513;
    'h03DF: mem_data <= 32'hB6CFF0EF;
    'h03E0: mem_data <= 32'h001027B7;
    'h03E1: mem_data <= 32'hCC078513;
    'h03E2: mem_data <= 32'hA60FF0EF;
    'h03E3: mem_data <= 32'h00304783;
    'h03E4: mem_data <= 32'h00078513;
    'h03E5: mem_data <= 32'hB54FF0EF;
    'h03E6: mem_data <= 32'h001027B7;
    'h03E7: mem_data <= 32'hAD878513;
    'h03E8: mem_data <= 32'hA48FF0EF;
    'h03E9: mem_data <= 32'h00000223;
    'h03EA: mem_data <= 32'h23C0006F;
    'h03EB: mem_data <= 32'h00204783;
    'h03EC: mem_data <= 32'h00379793;
    'h03ED: mem_data <= 32'h0087F793;
    'h03EE: mem_data <= 32'h0D07E713;
    'h03EF: mem_data <= 32'h00304783;
    'h03F0: mem_data <= 32'h00279793;
    'h03F1: mem_data <= 32'h0047F793;
    'h03F2: mem_data <= 32'h00F76733;
    'h03F3: mem_data <= 32'h00404783;
    'h03F4: mem_data <= 32'h0037F793;
    'h03F5: mem_data <= 32'h00F76733;
    'h03F6: mem_data <= 32'h050007B7;
    'h03F7: mem_data <= 32'h00E7A023;
    'h03F8: mem_data <= 32'h050007B7;
    'h03F9: mem_data <= 32'h40078793;
    'h03FA: mem_data <= 32'hFCF44703;
    'h03FB: mem_data <= 32'h00E7A023;
    'h03FC: mem_data <= 32'h050007B7;
    'h03FD: mem_data <= 32'h30078793;
    'h03FE: mem_data <= 32'h0007A023;
    'h03FF: mem_data <= 32'h001027B7;
    'h0400: mem_data <= 32'hC6078513;
    'h0401: mem_data <= 32'h9E4FF0EF;
    'h0402: mem_data <= 32'h000002A3;
    'h0403: mem_data <= 32'h0E00006F;
    'h0404: mem_data <= 32'h00204783;
    'h0405: mem_data <= 32'h00779793;
    'h0406: mem_data <= 32'h01879713;
    'h0407: mem_data <= 32'h41875713;
    'h0408: mem_data <= 32'h00304783;
    'h0409: mem_data <= 32'h00679793;
    'h040A: mem_data <= 32'h01879793;
    'h040B: mem_data <= 32'h4187D793;
    'h040C: mem_data <= 32'h0407F793;
    'h040D: mem_data <= 32'h01879793;
    'h040E: mem_data <= 32'h4187D793;
    'h040F: mem_data <= 32'h00F767B3;
    'h0410: mem_data <= 32'h01879713;
    'h0411: mem_data <= 32'h41875713;
    'h0412: mem_data <= 32'h00404783;
    'h0413: mem_data <= 32'h00479793;
    'h0414: mem_data <= 32'h01879793;
    'h0415: mem_data <= 32'h4187D793;
    'h0416: mem_data <= 32'h0307F793;
    'h0417: mem_data <= 32'h01879793;
    'h0418: mem_data <= 32'h4187D793;
    'h0419: mem_data <= 32'h00F767B3;
    'h041A: mem_data <= 32'h01879713;
    'h041B: mem_data <= 32'h41875713;
    'h041C: mem_data <= 32'h00504783;
    'h041D: mem_data <= 32'h01879793;
    'h041E: mem_data <= 32'h4187D793;
    'h041F: mem_data <= 32'h00F7F793;
    'h0420: mem_data <= 32'h01879793;
    'h0421: mem_data <= 32'h4187D793;
    'h0422: mem_data <= 32'h00F767B3;
    'h0423: mem_data <= 32'h01879793;
    'h0424: mem_data <= 32'h4187D793;
    'h0425: mem_data <= 32'h0FF7F713;
    'h0426: mem_data <= 32'h00E00423;
    'h0427: mem_data <= 32'h00804783;
    'h0428: mem_data <= 32'h00078513;
    'h0429: mem_data <= 32'hE19FF0EF;
    'h042A: mem_data <= 32'h00504783;
    'h042B: mem_data <= 32'h00078693;
    'h042C: mem_data <= 32'h00804703;
    'h042D: mem_data <= 32'hFF068793;
    'h042E: mem_data <= 32'h008787B3;
    'h042F: mem_data <= 32'hFEE78A23;
    'h0430: mem_data <= 32'h00804783;
    'h0431: mem_data <= 32'h00200593;
    'h0432: mem_data <= 32'h00078513;
    'h0433: mem_data <= 32'h970FF0EF;
    'h0434: mem_data <= 32'h001027B7;
    'h0435: mem_data <= 32'hC6C78513;
    'h0436: mem_data <= 32'h910FF0EF;
    'h0437: mem_data <= 32'h00504783;
    'h0438: mem_data <= 32'h00178793;
    'h0439: mem_data <= 32'h0FF7F713;
    'h043A: mem_data <= 32'h00E002A3;
    'h043B: mem_data <= 32'h00504703;
    'h043C: mem_data <= 32'h00700793;
    'h043D: mem_data <= 32'hF0E7FEE3;
    'h043E: mem_data <= 32'h001027B7;
    'h043F: mem_data <= 32'hC7078513;
    'h0440: mem_data <= 32'h8E8FF0EF;
    'h0441: mem_data <= 32'h000002A3;
    'h0442: mem_data <= 32'h06C0006F;
    'h0443: mem_data <= 32'h00504783;
    'h0444: mem_data <= 32'hFFF7C793;
    'h0445: mem_data <= 32'h0FF7F793;
    'h0446: mem_data <= 32'h00078513;
    'h0447: mem_data <= 32'hDA1FF0EF;
    'h0448: mem_data <= 32'h050107B7;
    'h0449: mem_data <= 32'h0007A783;
    'h044A: mem_data <= 32'h0FF7F713;
    'h044B: mem_data <= 32'h00E003A3;
    'h044C: mem_data <= 32'h00504783;
    'h044D: mem_data <= 32'h00078693;
    'h044E: mem_data <= 32'h00704703;
    'h044F: mem_data <= 32'hFF068793;
    'h0450: mem_data <= 32'h008787B3;
    'h0451: mem_data <= 32'hFEE78623;
    'h0452: mem_data <= 32'h00704783;
    'h0453: mem_data <= 32'h00200593;
    'h0454: mem_data <= 32'h00078513;
    'h0455: mem_data <= 32'h8E8FF0EF;
    'h0456: mem_data <= 32'h001027B7;
    'h0457: mem_data <= 32'hC6C78513;
    'h0458: mem_data <= 32'h888FF0EF;
    'h0459: mem_data <= 32'h00504783;
    'h045A: mem_data <= 32'h00178793;
    'h045B: mem_data <= 32'h0FF7F713;
    'h045C: mem_data <= 32'h00E002A3;
    'h045D: mem_data <= 32'h00504703;
    'h045E: mem_data <= 32'h00700793;
    'h045F: mem_data <= 32'hF8E7F8E3;
    'h0460: mem_data <= 32'h000002A3;
    'h0461: mem_data <= 32'h0440006F;
    'h0462: mem_data <= 32'h00504783;
    'h0463: mem_data <= 32'hFF078793;
    'h0464: mem_data <= 32'h008787B3;
    'h0465: mem_data <= 32'hFF47C703;
    'h0466: mem_data <= 32'h00504783;
    'h0467: mem_data <= 32'hFF078793;
    'h0468: mem_data <= 32'h008787B3;
    'h0469: mem_data <= 32'hFEC7C783;
    'h046A: mem_data <= 32'h00F71863;
    'h046B: mem_data <= 32'hFEF44783;
    'h046C: mem_data <= 32'h00178793;
    'h046D: mem_data <= 32'hFEF407A3;
    'h046E: mem_data <= 32'h00504783;
    'h046F: mem_data <= 32'h00178793;
    'h0470: mem_data <= 32'h0FF7F713;
    'h0471: mem_data <= 32'h00E002A3;
    'h0472: mem_data <= 32'h00504703;
    'h0473: mem_data <= 32'h00700793;
    'h0474: mem_data <= 32'hFAE7FCE3;
    'h0475: mem_data <= 32'h00404783;
    'h0476: mem_data <= 32'h00178793;
    'h0477: mem_data <= 32'h0FF7F713;
    'h0478: mem_data <= 32'h00E00223;
    'h0479: mem_data <= 32'h00404703;
    'h047A: mem_data <= 32'h00300793;
    'h047B: mem_data <= 32'hDCE7F0E3;
    'h047C: mem_data <= 32'h00304783;
    'h047D: mem_data <= 32'h00178793;
    'h047E: mem_data <= 32'h0FF7F713;
    'h047F: mem_data <= 32'h00E001A3;
    'h0480: mem_data <= 32'h00304703;
    'h0481: mem_data <= 32'h00100793;
    'h0482: mem_data <= 32'hD4E7F8E3;
    'h0483: mem_data <= 32'h00204783;
    'h0484: mem_data <= 32'h00178793;
    'h0485: mem_data <= 32'h0FF7F713;
    'h0486: mem_data <= 32'h00E00123;
    'h0487: mem_data <= 32'h00204703;
    'h0488: mem_data <= 32'h00100793;
    'h0489: mem_data <= 32'hD2E7F6E3;
    'h048A: mem_data <= 32'hFEF44703;
    'h048B: mem_data <= 32'h08000793;
    'h048C: mem_data <= 32'h00F71A63;
    'h048D: mem_data <= 32'h001027B7;
    'h048E: mem_data <= 32'hCCC78513;
    'h048F: mem_data <= 32'hFADFE0EF;
    'h0490: mem_data <= 32'h0100006F;
    'h0491: mem_data <= 32'h001027B7;
    'h0492: mem_data <= 32'hCE078513;
    'h0493: mem_data <= 32'hF9DFE0EF;
    'h0494: mem_data <= 32'h050007B7;
    'h0495: mem_data <= 32'h30078793;
    'h0496: mem_data <= 32'h00100713;
    'h0497: mem_data <= 32'h00E7A023;
    'h0498: mem_data <= 32'h050007B7;
    'h0499: mem_data <= 32'h01000713;
    'h049A: mem_data <= 32'h00E7A023;
    'h049B: mem_data <= 32'h00000013;
    'h049C: mem_data <= 32'h03C12083;
    'h049D: mem_data <= 32'h03812403;
    'h049E: mem_data <= 32'h04010113;
    'h049F: mem_data <= 32'h00008067;
    'h04A0: mem_data <= 32'hFF010113;
    'h04A1: mem_data <= 32'h00112623;
    'h04A2: mem_data <= 32'h00812423;
    'h04A3: mem_data <= 32'h01010413;
    'h04A4: mem_data <= 32'h001027B7;
    'h04A5: mem_data <= 32'hCF878513;
    'h04A6: mem_data <= 32'hF51FE0EF;
    'h04A7: mem_data <= 32'h00000013;
    'h04A8: mem_data <= 32'h00C12083;
    'h04A9: mem_data <= 32'h00812403;
    'h04AA: mem_data <= 32'h01010113;
    'h04AB: mem_data <= 32'h00008067;
    'h04AC: mem_data <= 32'hFE010113;
    'h04AD: mem_data <= 32'h00112E23;
    'h04AE: mem_data <= 32'h00812C23;
    'h04AF: mem_data <= 32'h02010413;
    'h04B0: mem_data <= 32'h00A00793;
    'h04B1: mem_data <= 32'hFEF42623;
    'h04B2: mem_data <= 32'h00000013;
    'h04B3: mem_data <= 32'hFEC42783;
    'h04B4: mem_data <= 32'h04F05C63;
    'h04B5: mem_data <= 32'h001027B7;
    'h04B6: mem_data <= 32'hD0478513;
    'h04B7: mem_data <= 32'hF0DFE0EF;
    'h04B8: mem_data <= 32'hB80FF0EF;
    'h04B9: mem_data <= 32'h00050793;
    'h04BA: mem_data <= 32'hFEF405A3;
    'h04BB: mem_data <= 32'hFEB44703;
    'h04BC: mem_data <= 32'h02000793;
    'h04BD: mem_data <= 32'h00E7FE63;
    'h04BE: mem_data <= 32'hFEB44703;
    'h04BF: mem_data <= 32'h07E00793;
    'h04C0: mem_data <= 32'h00E7E863;
    'h04C1: mem_data <= 32'hFEB44783;
    'h04C2: mem_data <= 32'h00078513;
    'h04C3: mem_data <= 32'hE8DFE0EF;
    'h04C4: mem_data <= 32'h001027B7;
    'h04C5: mem_data <= 32'hAD878513;
    'h04C6: mem_data <= 32'hED1FE0EF;
    'h04C7: mem_data <= 32'h00000013;
    'h04C8: mem_data <= 32'hF61FF0EF;
    'h04C9: mem_data <= 32'h0080006F;
    'h04CA: mem_data <= 32'h00000013;
    'h04CB: mem_data <= 32'h00000013;
    'h04CC: mem_data <= 32'h01C12083;
    'h04CD: mem_data <= 32'h01812403;
    'h04CE: mem_data <= 32'h02010113;
    'h04CF: mem_data <= 32'h00008067;
    'h04D0: mem_data <= 32'hFE010113;
    'h04D1: mem_data <= 32'h00112E23;
    'h04D2: mem_data <= 32'h00812C23;
    'h04D3: mem_data <= 32'h02010413;
    'h04D4: mem_data <= 32'h00A00793;
    'h04D5: mem_data <= 32'hFEF42623;
    'h04D6: mem_data <= 32'h0740006F;
    'h04D7: mem_data <= 32'h001027B7;
    'h04D8: mem_data <= 32'hD2478513;
    'h04D9: mem_data <= 32'hE85FE0EF;
    'h04DA: mem_data <= 32'hAF8FF0EF;
    'h04DB: mem_data <= 32'h00050793;
    'h04DC: mem_data <= 32'hFEF405A3;
    'h04DD: mem_data <= 32'hFEB44703;
    'h04DE: mem_data <= 32'h02000793;
    'h04DF: mem_data <= 32'h00E7FE63;
    'h04E0: mem_data <= 32'hFEB44703;
    'h04E1: mem_data <= 32'h07E00793;
    'h04E2: mem_data <= 32'h00E7E863;
    'h04E3: mem_data <= 32'hFEB44783;
    'h04E4: mem_data <= 32'h00078513;
    'h04E5: mem_data <= 32'hE05FE0EF;
    'h04E6: mem_data <= 32'h001027B7;
    'h04E7: mem_data <= 32'hAD878513;
    'h04E8: mem_data <= 32'hE49FE0EF;
    'h04E9: mem_data <= 32'hFEB44703;
    'h04EA: mem_data <= 32'h00D00793;
    'h04EB: mem_data <= 32'h00F71863;
    'h04EC: mem_data <= 32'h00000013;
    'h04ED: mem_data <= 32'hECDFF0EF;
    'h04EE: mem_data <= 32'h0200006F;
    'h04EF: mem_data <= 32'h00000013;
    'h04F0: mem_data <= 32'hFEC42783;
    'h04F1: mem_data <= 32'hFFF78793;
    'h04F2: mem_data <= 32'hFEF42623;
    'h04F3: mem_data <= 32'hFEC42783;
    'h04F4: mem_data <= 32'hF8F046E3;
    'h04F5: mem_data <= 32'h00000013;
    'h04F6: mem_data <= 32'h00000013;
    'h04F7: mem_data <= 32'h01C12083;
    'h04F8: mem_data <= 32'h01812403;
    'h04F9: mem_data <= 32'h02010113;
    'h04FA: mem_data <= 32'h00008067;
    'h04FB: mem_data <= 32'hFF010113;
    'h04FC: mem_data <= 32'h00112623;
    'h04FD: mem_data <= 32'h00812423;
    'h04FE: mem_data <= 32'h01010413;
    'h04FF: mem_data <= 32'h001027B7;
    'h0500: mem_data <= 32'hD4078513;
    'h0501: mem_data <= 32'hDE5FE0EF;
    'h0502: mem_data <= 32'h00000013;
    'h0503: mem_data <= 32'h00C12083;
    'h0504: mem_data <= 32'h00812403;
    'h0505: mem_data <= 32'h01010113;
    'h0506: mem_data <= 32'h00008067;
    'h0507: mem_data <= 32'hFF010113;
    'h0508: mem_data <= 32'h00112623;
    'h0509: mem_data <= 32'h00812423;
    'h050A: mem_data <= 32'h01010413;
    'h050B: mem_data <= 32'h030007B7;
    'h050C: mem_data <= 32'h00100713;
    'h050D: mem_data <= 32'h00E7A023;
    'h050E: mem_data <= 32'h001027B7;
    'h050F: mem_data <= 32'hF4078513;
    'h0510: mem_data <= 32'hDA9FE0EF;
    'h0511: mem_data <= 32'h00000013;
    'h0512: mem_data <= 32'h00C12083;
    'h0513: mem_data <= 32'h00812403;
    'h0514: mem_data <= 32'h01010113;
    'h0515: mem_data <= 32'h00008067;
    'h0516: mem_data <= 32'hFF010113;
    'h0517: mem_data <= 32'h00112623;
    'h0518: mem_data <= 32'h00812423;
    'h0519: mem_data <= 32'h01010413;
    'h051A: mem_data <= 32'h030007B7;
    'h051B: mem_data <= 32'h00200713;
    'h051C: mem_data <= 32'h00E7A023;
    'h051D: mem_data <= 32'h001037B7;
    'h051E: mem_data <= 32'h88C78513;
    'h051F: mem_data <= 32'hD6DFE0EF;
    'h0520: mem_data <= 32'h00000013;
    'h0521: mem_data <= 32'h00C12083;
    'h0522: mem_data <= 32'h00812403;
    'h0523: mem_data <= 32'h01010113;
    'h0524: mem_data <= 32'h00008067;
    'h0525: mem_data <= 32'hFE010113;
    'h0526: mem_data <= 32'h00112E23;
    'h0527: mem_data <= 32'h00812C23;
    'h0528: mem_data <= 32'h02010413;
    'h0529: mem_data <= 32'h030007B7;
    'h052A: mem_data <= 32'h0FF00713;
    'h052B: mem_data <= 32'h00E7A023;
    'h052C: mem_data <= 32'hF3DFF0EF;
    'h052D: mem_data <= 32'h001037B7;
    'h052E: mem_data <= 32'hAC078513;
    'h052F: mem_data <= 32'hD2DFE0EF;
    'h0530: mem_data <= 32'h00A00793;
    'h0531: mem_data <= 32'hFEF42623;
    'h0532: mem_data <= 32'h0D00006F;
    'h0533: mem_data <= 32'h001037B7;
    'h0534: mem_data <= 32'hB2C78513;
    'h0535: mem_data <= 32'hD15FE0EF;
    'h0536: mem_data <= 32'h988FF0EF;
    'h0537: mem_data <= 32'h00050793;
    'h0538: mem_data <= 32'hFEF405A3;
    'h0539: mem_data <= 32'hFEB44703;
    'h053A: mem_data <= 32'h02000793;
    'h053B: mem_data <= 32'h00E7FE63;
    'h053C: mem_data <= 32'hFEB44703;
    'h053D: mem_data <= 32'h07E00793;
    'h053E: mem_data <= 32'h00E7E863;
    'h053F: mem_data <= 32'hFEB44783;
    'h0540: mem_data <= 32'h00078513;
    'h0541: mem_data <= 32'hC95FE0EF;
    'h0542: mem_data <= 32'h001027B7;
    'h0543: mem_data <= 32'hAD878513;
    'h0544: mem_data <= 32'hCD9FE0EF;
    'h0545: mem_data <= 32'hFEB44783;
    'h0546: mem_data <= 32'hFCF78793;
    'h0547: mem_data <= 32'h00400713;
    'h0548: mem_data <= 32'h06F76463;
    'h0549: mem_data <= 32'h00279713;
    'h054A: mem_data <= 32'h001037B7;
    'h054B: mem_data <= 32'hB3C78793;
    'h054C: mem_data <= 32'h00F707B3;
    'h054D: mem_data <= 32'h0007A783;
    'h054E: mem_data <= 32'h00078067;
    'h054F: mem_data <= 32'hD45FF0EF;
    'h0550: mem_data <= 32'hEDDFF0EF;
    'h0551: mem_data <= 32'hD6DFF0EF;
    'h0552: mem_data <= 32'h0380006F;
    'h0553: mem_data <= 32'hD35FF0EF;
    'h0554: mem_data <= 32'hF09FF0EF;
    'h0555: mem_data <= 32'hD5DFF0EF;
    'h0556: mem_data <= 32'h0280006F;
    'h0557: mem_data <= 32'hD25FF0EF;
    'h0558: mem_data <= 32'h058000EF;
    'h0559: mem_data <= 32'h01C0006F;
    'h055A: mem_data <= 32'hD19FF0EF;
    'h055B: mem_data <= 32'h158000EF;
    'h055C: mem_data <= 32'h0100006F;
    'h055D: mem_data <= 32'hD0DFF0EF;
    'h055E: mem_data <= 32'h264000EF;
    'h055F: mem_data <= 32'h00000013;
    'h0560: mem_data <= 32'hD01FF0EF;
    'h0561: mem_data <= 32'h0200006F;
    'h0562: mem_data <= 32'h00000013;
    'h0563: mem_data <= 32'hFEC42783;
    'h0564: mem_data <= 32'hFFF78793;
    'h0565: mem_data <= 32'hFEF42623;
    'h0566: mem_data <= 32'hFEC42783;
    'h0567: mem_data <= 32'hF2F048E3;
    'h0568: mem_data <= 32'h00000013;
    'h0569: mem_data <= 32'h00000013;
    'h056A: mem_data <= 32'h01C12083;
    'h056B: mem_data <= 32'h01812403;
    'h056C: mem_data <= 32'h02010113;
    'h056D: mem_data <= 32'h00008067;
    'h056E: mem_data <= 32'hFE010113;
    'h056F: mem_data <= 32'h00112E23;
    'h0570: mem_data <= 32'h00812C23;
    'h0571: mem_data <= 32'h02010413;
    'h0572: mem_data <= 32'h030007B7;
    'h0573: mem_data <= 32'h00300713;
    'h0574: mem_data <= 32'h00E7A023;
    'h0575: mem_data <= 32'hE19FF0EF;
    'h0576: mem_data <= 32'h001037B7;
    'h0577: mem_data <= 32'hB5078513;
    'h0578: mem_data <= 32'hC09FE0EF;
    'h0579: mem_data <= 32'h00A00793;
    'h057A: mem_data <= 32'hFEF42623;
    'h057B: mem_data <= 32'h0B80006F;
    'h057C: mem_data <= 32'h001037B7;
    'h057D: mem_data <= 32'hBB478513;
    'h057E: mem_data <= 32'hBF1FE0EF;
    'h057F: mem_data <= 32'h864FF0EF;
    'h0580: mem_data <= 32'h00050793;
    'h0581: mem_data <= 32'hFEF405A3;
    'h0582: mem_data <= 32'hFEB44703;
    'h0583: mem_data <= 32'h02000793;
    'h0584: mem_data <= 32'h00E7FE63;
    'h0585: mem_data <= 32'hFEB44703;
    'h0586: mem_data <= 32'h07E00793;
    'h0587: mem_data <= 32'h00E7E863;
    'h0588: mem_data <= 32'hFEB44783;
    'h0589: mem_data <= 32'h00078513;
    'h058A: mem_data <= 32'hB71FE0EF;
    'h058B: mem_data <= 32'h001027B7;
    'h058C: mem_data <= 32'hAD878513;
    'h058D: mem_data <= 32'hBB5FE0EF;
    'h058E: mem_data <= 32'hFEB44783;
    'h058F: mem_data <= 32'h07200713;
    'h0590: mem_data <= 32'h02E78E63;
    'h0591: mem_data <= 32'h07200713;
    'h0592: mem_data <= 32'h04F74663;
    'h0593: mem_data <= 32'h03100713;
    'h0594: mem_data <= 32'h00E78863;
    'h0595: mem_data <= 32'h03200713;
    'h0596: mem_data <= 32'h00E78A63;
    'h0597: mem_data <= 32'h0380006F;
    'h0598: mem_data <= 32'hC21FF0EF;
    'h0599: mem_data <= 32'h8A0FF0EF;
    'h059A: mem_data <= 32'h0240006F;
    'h059B: mem_data <= 32'hC15FF0EF;
    'h059C: mem_data <= 32'hA2CFF0EF;
    'h059D: mem_data <= 32'hC3DFF0EF;
    'h059E: mem_data <= 32'h0140006F;
    'h059F: mem_data <= 32'hC05FF0EF;
    'h05A0: mem_data <= 32'hE15FF0EF;
    'h05A1: mem_data <= 32'hC2DFF0EF;
    'h05A2: mem_data <= 32'h00000013;
    'h05A3: mem_data <= 32'hBF5FF0EF;
    'h05A4: mem_data <= 32'h0200006F;
    'h05A5: mem_data <= 32'h00000013;
    'h05A6: mem_data <= 32'hFEC42783;
    'h05A7: mem_data <= 32'hFFF78793;
    'h05A8: mem_data <= 32'hFEF42623;
    'h05A9: mem_data <= 32'hFEC42783;
    'h05AA: mem_data <= 32'hF4F044E3;
    'h05AB: mem_data <= 32'h00000013;
    'h05AC: mem_data <= 32'h00000013;
    'h05AD: mem_data <= 32'h01C12083;
    'h05AE: mem_data <= 32'h01812403;
    'h05AF: mem_data <= 32'h02010113;
    'h05B0: mem_data <= 32'h00008067;
    'h05B1: mem_data <= 32'hFE010113;
    'h05B2: mem_data <= 32'h00112E23;
    'h05B3: mem_data <= 32'h00812C23;
    'h05B4: mem_data <= 32'h02010413;
    'h05B5: mem_data <= 32'h030007B7;
    'h05B6: mem_data <= 32'h00400713;
    'h05B7: mem_data <= 32'h00E7A023;
    'h05B8: mem_data <= 32'hD0DFF0EF;
    'h05B9: mem_data <= 32'h001037B7;
    'h05BA: mem_data <= 32'hBC478513;
    'h05BB: mem_data <= 32'hAFDFE0EF;
    'h05BC: mem_data <= 32'h00A00793;
    'h05BD: mem_data <= 32'hFEF42623;
    'h05BE: mem_data <= 32'h0C40006F;
    'h05BF: mem_data <= 32'h001037B7;
    'h05C0: mem_data <= 32'hBB478513;
    'h05C1: mem_data <= 32'hAE5FE0EF;
    'h05C2: mem_data <= 32'hF59FE0EF;
    'h05C3: mem_data <= 32'h00050793;
    'h05C4: mem_data <= 32'hFEF405A3;
    'h05C5: mem_data <= 32'hFEB44703;
    'h05C6: mem_data <= 32'h02000793;
    'h05C7: mem_data <= 32'h00E7FE63;
    'h05C8: mem_data <= 32'hFEB44703;
    'h05C9: mem_data <= 32'h07E00793;
    'h05CA: mem_data <= 32'h00E7E863;
    'h05CB: mem_data <= 32'hFEB44783;
    'h05CC: mem_data <= 32'h00078513;
    'h05CD: mem_data <= 32'hA65FE0EF;
    'h05CE: mem_data <= 32'h001027B7;
    'h05CF: mem_data <= 32'hAD878513;
    'h05D0: mem_data <= 32'hAA9FE0EF;
    'h05D1: mem_data <= 32'hFEB44783;
    'h05D2: mem_data <= 32'h07200713;
    'h05D3: mem_data <= 32'h04E78463;
    'h05D4: mem_data <= 32'h07200713;
    'h05D5: mem_data <= 32'h04F74C63;
    'h05D6: mem_data <= 32'h03100713;
    'h05D7: mem_data <= 32'h00E78863;
    'h05D8: mem_data <= 32'h03200713;
    'h05D9: mem_data <= 32'h00E78E63;
    'h05DA: mem_data <= 32'h0440006F;
    'h05DB: mem_data <= 32'hB15FF0EF;
    'h05DC: mem_data <= 32'h07D00513;
    'h05DD: mem_data <= 32'hC68FF0EF;
    'h05DE: mem_data <= 32'hB39FF0EF;
    'h05DF: mem_data <= 32'h0280006F;
    'h05E0: mem_data <= 32'hB01FF0EF;
    'h05E1: mem_data <= 32'h01F00513;
    'h05E2: mem_data <= 32'hC54FF0EF;
    'h05E3: mem_data <= 32'hB25FF0EF;
    'h05E4: mem_data <= 32'h0140006F;
    'h05E5: mem_data <= 32'hAEDFF0EF;
    'h05E6: mem_data <= 32'hCFDFF0EF;
    'h05E7: mem_data <= 32'hB15FF0EF;
    'h05E8: mem_data <= 32'h00000013;
    'h05E9: mem_data <= 32'hADDFF0EF;
    'h05EA: mem_data <= 32'h0200006F;
    'h05EB: mem_data <= 32'h00000013;
    'h05EC: mem_data <= 32'hFEC42783;
    'h05ED: mem_data <= 32'hFFF78793;
    'h05EE: mem_data <= 32'hFEF42623;
    'h05EF: mem_data <= 32'hFEC42783;
    'h05F0: mem_data <= 32'hF2F04EE3;
    'h05F1: mem_data <= 32'h00000013;
    'h05F2: mem_data <= 32'h00000013;
    'h05F3: mem_data <= 32'h01C12083;
    'h05F4: mem_data <= 32'h01812403;
    'h05F5: mem_data <= 32'h02010113;
    'h05F6: mem_data <= 32'h00008067;
    'h05F7: mem_data <= 32'hFE010113;
    'h05F8: mem_data <= 32'h00112E23;
    'h05F9: mem_data <= 32'h00812C23;
    'h05FA: mem_data <= 32'h02010413;
    'h05FB: mem_data <= 32'h030007B7;
    'h05FC: mem_data <= 32'h00500713;
    'h05FD: mem_data <= 32'h00E7A023;
    'h05FE: mem_data <= 32'hBF5FF0EF;
    'h05FF: mem_data <= 32'h001037B7;
    'h0600: mem_data <= 32'hC3078513;
    'h0601: mem_data <= 32'h9E5FE0EF;
    'h0602: mem_data <= 32'h00A00793;
    'h0603: mem_data <= 32'hFEF42623;
    'h0604: mem_data <= 32'h10C0006F;
    'h0605: mem_data <= 32'h001037B7;
    'h0606: mem_data <= 32'hCE878513;
    'h0607: mem_data <= 32'h9CDFE0EF;
    'h0608: mem_data <= 32'hE41FE0EF;
    'h0609: mem_data <= 32'h00050793;
    'h060A: mem_data <= 32'hFEF405A3;
    'h060B: mem_data <= 32'hFEB44703;
    'h060C: mem_data <= 32'h02000793;
    'h060D: mem_data <= 32'h00E7FE63;
    'h060E: mem_data <= 32'hFEB44703;
    'h060F: mem_data <= 32'h07E00793;
    'h0610: mem_data <= 32'h00E7E863;
    'h0611: mem_data <= 32'hFEB44783;
    'h0612: mem_data <= 32'h00078513;
    'h0613: mem_data <= 32'h94DFE0EF;
    'h0614: mem_data <= 32'h001027B7;
    'h0615: mem_data <= 32'hAD878513;
    'h0616: mem_data <= 32'h991FE0EF;
    'h0617: mem_data <= 32'hFEB44783;
    'h0618: mem_data <= 32'h07200713;
    'h0619: mem_data <= 32'h08E78863;
    'h061A: mem_data <= 32'h07200713;
    'h061B: mem_data <= 32'h0AF74063;
    'h061C: mem_data <= 32'h03400713;
    'h061D: mem_data <= 32'h06E78663;
    'h061E: mem_data <= 32'h03400713;
    'h061F: mem_data <= 32'h08F74863;
    'h0620: mem_data <= 32'h03300713;
    'h0621: mem_data <= 32'h04E78463;
    'h0622: mem_data <= 32'h03300713;
    'h0623: mem_data <= 32'h08F74063;
    'h0624: mem_data <= 32'h03100713;
    'h0625: mem_data <= 32'h00E78863;
    'h0626: mem_data <= 32'h03200713;
    'h0627: mem_data <= 32'h00E78E63;
    'h0628: mem_data <= 32'h06C0006F;
    'h0629: mem_data <= 32'h9DDFF0EF;
    'h062A: mem_data <= 32'h0D800513;
    'h062B: mem_data <= 32'hE50FF0EF;
    'h062C: mem_data <= 32'hA01FF0EF;
    'h062D: mem_data <= 32'h0500006F;
    'h062E: mem_data <= 32'h9C9FF0EF;
    'h062F: mem_data <= 32'h06B00513;
    'h0630: mem_data <= 32'hE3CFF0EF;
    'h0631: mem_data <= 32'h9EDFF0EF;
    'h0632: mem_data <= 32'h03C0006F;
    'h0633: mem_data <= 32'h9B5FF0EF;
    'h0634: mem_data <= 32'h03500513;
    'h0635: mem_data <= 32'hE28FF0EF;
    'h0636: mem_data <= 32'h9D9FF0EF;
    'h0637: mem_data <= 32'h0280006F;
    'h0638: mem_data <= 32'h9A1FF0EF;
    'h0639: mem_data <= 32'h01A00513;
    'h063A: mem_data <= 32'hE14FF0EF;
    'h063B: mem_data <= 32'h9C5FF0EF;
    'h063C: mem_data <= 32'h0140006F;
    'h063D: mem_data <= 32'h98DFF0EF;
    'h063E: mem_data <= 32'hB9DFF0EF;
    'h063F: mem_data <= 32'h9B5FF0EF;
    'h0640: mem_data <= 32'h00000013;
    'h0641: mem_data <= 32'h97DFF0EF;
    'h0642: mem_data <= 32'h0200006F;
    'h0643: mem_data <= 32'h00000013;
    'h0644: mem_data <= 32'hFEC42783;
    'h0645: mem_data <= 32'hFFF78793;
    'h0646: mem_data <= 32'hFEF42623;
    'h0647: mem_data <= 32'hFEC42783;
    'h0648: mem_data <= 32'hEEF04AE3;
    'h0649: mem_data <= 32'h00000013;
    'h064A: mem_data <= 32'h00000013;
    'h064B: mem_data <= 32'h01C12083;
    'h064C: mem_data <= 32'h01812403;
    'h064D: mem_data <= 32'h02010113;
    'h064E: mem_data <= 32'h00008067;
    'h064F: mem_data <= 32'hFF010113;
    'h0650: mem_data <= 32'h00112623;
    'h0651: mem_data <= 32'h00812423;
    'h0652: mem_data <= 32'h01010413;
    'h0653: mem_data <= 32'h020007B7;
    'h0654: mem_data <= 32'h00478793;
    'h0655: mem_data <= 32'h1B200713;
    'h0656: mem_data <= 32'h00E7A023;
    'h0657: mem_data <= 32'h030007B7;
    'h0658: mem_data <= 32'h01800713;
    'h0659: mem_data <= 32'h00E7A023;
    'h065A: mem_data <= 32'h0C800513;
    'h065B: mem_data <= 32'hD25FE0EF;
    'h065C: mem_data <= 32'h911FF0EF;
    'h065D: mem_data <= 32'h030007B7;
    'h065E: mem_data <= 32'h0FF00713;
    'h065F: mem_data <= 32'h00E7A023;
    'h0660: mem_data <= 32'h001037B7;
    'h0661: mem_data <= 32'hCFC78513;
    'h0662: mem_data <= 32'h861FE0EF;
    'h0663: mem_data <= 32'h030007B7;
    'h0664: mem_data <= 32'h07F00713;
    'h0665: mem_data <= 32'h00E7A023;
    'h0666: mem_data <= 32'h001037B7;
    'h0667: mem_data <= 32'hD0478513;
    'h0668: mem_data <= 32'h849FE0EF;
    'h0669: mem_data <= 32'h00100513;
    'h066A: mem_data <= 32'hCE9FE0EF;
    'h066B: mem_data <= 32'h030007B7;
    'h066C: mem_data <= 32'h03F00713;
    'h066D: mem_data <= 32'h00E7A023;
    'h066E: mem_data <= 32'h001037B7;
    'h066F: mem_data <= 32'hD0478513;
    'h0670: mem_data <= 32'h829FE0EF;
    'h0671: mem_data <= 32'h00100513;
    'h0672: mem_data <= 32'hCC9FE0EF;
    'h0673: mem_data <= 32'h030007B7;
    'h0674: mem_data <= 32'h01F00713;
    'h0675: mem_data <= 32'h00E7A023;
    'h0676: mem_data <= 32'h001037B7;
    'h0677: mem_data <= 32'hD0478513;
    'h0678: mem_data <= 32'h809FE0EF;
    'h0679: mem_data <= 32'h00100513;
    'h067A: mem_data <= 32'hCA9FE0EF;
    'h067B: mem_data <= 32'h030007B7;
    'h067C: mem_data <= 32'h00F00713;
    'h067D: mem_data <= 32'h00E7A023;
    'h067E: mem_data <= 32'h001037B7;
    'h067F: mem_data <= 32'hD0478513;
    'h0680: mem_data <= 32'hFE8FE0EF;
    'h0681: mem_data <= 32'h00100513;
    'h0682: mem_data <= 32'hC89FE0EF;
    'h0683: mem_data <= 32'h030007B7;
    'h0684: mem_data <= 32'h00700713;
    'h0685: mem_data <= 32'h00E7A023;
    'h0686: mem_data <= 32'h001037B7;
    'h0687: mem_data <= 32'hD0478513;
    'h0688: mem_data <= 32'hFC8FE0EF;
    'h0689: mem_data <= 32'h00100513;
    'h068A: mem_data <= 32'hC69FE0EF;
    'h068B: mem_data <= 32'h030007B7;
    'h068C: mem_data <= 32'h00300713;
    'h068D: mem_data <= 32'h00E7A023;
    'h068E: mem_data <= 32'h001037B7;
    'h068F: mem_data <= 32'hD0478513;
    'h0690: mem_data <= 32'hFA8FE0EF;
    'h0691: mem_data <= 32'h00100513;
    'h0692: mem_data <= 32'hC49FE0EF;
    'h0693: mem_data <= 32'h030007B7;
    'h0694: mem_data <= 32'h00100713;
    'h0695: mem_data <= 32'h00E7A023;
    'h0696: mem_data <= 32'h001037B7;
    'h0697: mem_data <= 32'hD0878513;
    'h0698: mem_data <= 32'hF88FE0EF;
    'h0699: mem_data <= 32'h00100513;
    'h069A: mem_data <= 32'hC29FE0EF;
    'h069B: mem_data <= 32'h030007B7;
    'h069C: mem_data <= 32'h0FF00713;
    'h069D: mem_data <= 32'h00E7A023;
    'h069E: mem_data <= 32'h8C9FF0EF;
    'h069F: mem_data <= 32'hA19FF0EF;
    'h06A0: mem_data <= 32'hFFDFF06F;
    'h06A1: mem_data <= 32'h33323130;
    'h06A2: mem_data <= 32'h37363534;
    'h06A3: mem_data <= 32'h42413938;
    'h06A4: mem_data <= 32'h46454443;
    'h06A5: mem_data <= 32'h00000000;
    'h06A6: mem_data <= 32'h30313D3E;
    'h06A7: mem_data <= 32'h00000030;
    'h06A8: mem_data <= 32'h73657250;
    'h06A9: mem_data <= 32'h20312073;
    'h06AA: mem_data <= 32'h38206F74;
    'h06AB: mem_data <= 32'h726F6620;
    'h06AC: mem_data <= 32'h72757420;
    'h06AD: mem_data <= 32'h6E6F206E;
    'h06AE: mem_data <= 32'h44454C20;
    'h06AF: mem_data <= 32'h20726F20;
    'h06B0: mem_data <= 32'h73657270;
    'h06B1: mem_data <= 32'h20522073;
    'h06B2: mem_data <= 32'h72206F74;
    'h06B3: mem_data <= 32'h72757465;
    'h06B4: mem_data <= 32'h2E2E2E6E;
    'h06B5: mem_data <= 32'h00000000;
    'h06B6: mem_data <= 32'h0000000A;
    'h06B7: mem_data <= 32'h00100798;
    'h06B8: mem_data <= 32'h001007B0;
    'h06B9: mem_data <= 32'h001007C8;
    'h06BA: mem_data <= 32'h001007E0;
    'h06BB: mem_data <= 32'h001007F8;
    'h06BC: mem_data <= 32'h00100810;
    'h06BD: mem_data <= 32'h00100828;
    'h06BE: mem_data <= 32'h00100840;
    'h06BF: mem_data <= 32'h0010086C;
    'h06C0: mem_data <= 32'h0010086C;
    'h06C1: mem_data <= 32'h0010086C;
    'h06C2: mem_data <= 32'h0010086C;
    'h06C3: mem_data <= 32'h0010086C;
    'h06C4: mem_data <= 32'h0010086C;
    'h06C5: mem_data <= 32'h0010086C;
    'h06C6: mem_data <= 32'h0010086C;
    'h06C7: mem_data <= 32'h0010086C;
    'h06C8: mem_data <= 32'h0010086C;
    'h06C9: mem_data <= 32'h0010086C;
    'h06CA: mem_data <= 32'h0010086C;
    'h06CB: mem_data <= 32'h0010086C;
    'h06CC: mem_data <= 32'h0010086C;
    'h06CD: mem_data <= 32'h0010086C;
    'h06CE: mem_data <= 32'h0010086C;
    'h06CF: mem_data <= 32'h0010086C;
    'h06D0: mem_data <= 32'h0010086C;
    'h06D1: mem_data <= 32'h0010086C;
    'h06D2: mem_data <= 32'h0010086C;
    'h06D3: mem_data <= 32'h0010086C;
    'h06D4: mem_data <= 32'h0010086C;
    'h06D5: mem_data <= 32'h0010086C;
    'h06D6: mem_data <= 32'h0010086C;
    'h06D7: mem_data <= 32'h0010086C;
    'h06D8: mem_data <= 32'h0010086C;
    'h06D9: mem_data <= 32'h0010086C;
    'h06DA: mem_data <= 32'h0010086C;
    'h06DB: mem_data <= 32'h0010086C;
    'h06DC: mem_data <= 32'h0010086C;
    'h06DD: mem_data <= 32'h0010086C;
    'h06DE: mem_data <= 32'h0010086C;
    'h06DF: mem_data <= 32'h0010086C;
    'h06E0: mem_data <= 32'h0010086C;
    'h06E1: mem_data <= 32'h0010086C;
    'h06E2: mem_data <= 32'h0010086C;
    'h06E3: mem_data <= 32'h0010086C;
    'h06E4: mem_data <= 32'h0010086C;
    'h06E5: mem_data <= 32'h0010086C;
    'h06E6: mem_data <= 32'h0010086C;
    'h06E7: mem_data <= 32'h0010086C;
    'h06E8: mem_data <= 32'h0010086C;
    'h06E9: mem_data <= 32'h0010086C;
    'h06EA: mem_data <= 32'h0010086C;
    'h06EB: mem_data <= 32'h0010086C;
    'h06EC: mem_data <= 32'h0010086C;
    'h06ED: mem_data <= 32'h0010086C;
    'h06EE: mem_data <= 32'h0010086C;
    'h06EF: mem_data <= 32'h0010086C;
    'h06F0: mem_data <= 32'h0010086C;
    'h06F1: mem_data <= 32'h0010086C;
    'h06F2: mem_data <= 32'h0010086C;
    'h06F3: mem_data <= 32'h0010086C;
    'h06F4: mem_data <= 32'h0010086C;
    'h06F5: mem_data <= 32'h0010086C;
    'h06F6: mem_data <= 32'h0010086C;
    'h06F7: mem_data <= 32'h0010086C;
    'h06F8: mem_data <= 32'h00100858;
    'h06F9: mem_data <= 32'h54545542;
    'h06FA: mem_data <= 32'h305F4E4F;
    'h06FB: mem_data <= 32'h00000020;
    'h06FC: mem_data <= 32'h0A46464F;
    'h06FD: mem_data <= 32'h00000000;
    'h06FE: mem_data <= 32'h000A4E4F;
    'h06FF: mem_data <= 32'h54545542;
    'h0700: mem_data <= 32'h315F4E4F;
    'h0701: mem_data <= 32'h00000020;
    'h0702: mem_data <= 32'h0A46464F;
    'h0703: mem_data <= 32'h0000000A;
    'h0704: mem_data <= 32'h0A0A4E4F;
    'h0705: mem_data <= 32'h00000000;
    'h0706: mem_data <= 32'h54495753;
    'h0707: mem_data <= 32'h305F4843;
    'h0708: mem_data <= 32'h00000020;
    'h0709: mem_data <= 32'h2D2D0A0A;
    'h070A: mem_data <= 32'h2D2D2D2D;
    'h070B: mem_data <= 32'h2D2D2D2D;
    'h070C: mem_data <= 32'h2D2D2D2D;
    'h070D: mem_data <= 32'h2D2D2D2D;
    'h070E: mem_data <= 32'h00000A2D;
    'h070F: mem_data <= 32'h54202020;
    'h0710: mem_data <= 32'h20545345;
    'h0711: mem_data <= 32'h00433249;
    'h0712: mem_data <= 32'h2D2D2D0A;
    'h0713: mem_data <= 32'h2D2D2D2D;
    'h0714: mem_data <= 32'h2D2D2D2D;
    'h0715: mem_data <= 32'h2D2D2D2D;
    'h0716: mem_data <= 32'h2D2D2D2D;
    'h0717: mem_data <= 32'h0000000A;
    'h0718: mem_data <= 32'h4952570A;
    'h0719: mem_data <= 32'h203A4554;
    'h071A: mem_data <= 32'h00000000;
    'h071B: mem_data <= 32'h00000020;
    'h071C: mem_data <= 32'h4145520A;
    'h071D: mem_data <= 32'h20203A44;
    'h071E: mem_data <= 32'h00000000;
    'h071F: mem_data <= 32'h65540A0A;
    'h0720: mem_data <= 32'h49207473;
    'h0721: mem_data <= 32'h70204332;
    'h0722: mem_data <= 32'h65737361;
    'h0723: mem_data <= 32'h000A2164;
    'h0724: mem_data <= 32'h65540A0A;
    'h0725: mem_data <= 32'h49207473;
    'h0726: mem_data <= 32'h6E204332;
    'h0727: mem_data <= 32'h7020746F;
    'h0728: mem_data <= 32'h65737361;
    'h0729: mem_data <= 32'h000A2164;
    'h072A: mem_data <= 32'h54202020;
    'h072B: mem_data <= 32'h20545345;
    'h072C: mem_data <= 32'h00495053;
    'h072D: mem_data <= 32'h50430A0A;
    'h072E: mem_data <= 32'h3D204C4F;
    'h072F: mem_data <= 32'h00000020;
    'h0730: mem_data <= 32'h20202020;
    'h0731: mem_data <= 32'h41485043;
    'h0732: mem_data <= 32'h00203D20;
    'h0733: mem_data <= 32'h65540A0A;
    'h0734: mem_data <= 32'h53207473;
    'h0735: mem_data <= 32'h70204950;
    'h0736: mem_data <= 32'h65737361;
    'h0737: mem_data <= 32'h000A2164;
    'h0738: mem_data <= 32'h65540A0A;
    'h0739: mem_data <= 32'h53207473;
    'h073A: mem_data <= 32'h6E204950;
    'h073B: mem_data <= 32'h7020746F;
    'h073C: mem_data <= 32'h65737361;
    'h073D: mem_data <= 32'h000A2164;
    'h073E: mem_data <= 32'h3B315B1B;
    'h073F: mem_data <= 32'h5B1B4831;
    'h0740: mem_data <= 32'h00004A32;
    'h0741: mem_data <= 32'h72500A0A;
    'h0742: mem_data <= 32'h20737365;
    'h0743: mem_data <= 32'h20796E61;
    'h0744: mem_data <= 32'h2079656B;
    'h0745: mem_data <= 32'h63206F74;
    'h0746: mem_data <= 32'h69746E6F;
    'h0747: mem_data <= 32'h2E65756E;
    'h0748: mem_data <= 32'h00002E2E;
    'h0749: mem_data <= 32'h73657250;
    'h074A: mem_data <= 32'h4E452073;
    'h074B: mem_data <= 32'h20524554;
    'h074C: mem_data <= 32'h63206F74;
    'h074D: mem_data <= 32'h69746E6F;
    'h074E: mem_data <= 32'h2E65756E;
    'h074F: mem_data <= 32'h00002E2E;
    'h0750: mem_data <= 32'h5F202020;
    'h0751: mem_data <= 32'h5F5F5F5F;
    'h0752: mem_data <= 32'h5F5F5F5F;
    'h0753: mem_data <= 32'h5F5F5F20;
    'h0754: mem_data <= 32'h5F5F5F5F;
    'h0755: mem_data <= 32'h5F5F2020;
    'h0756: mem_data <= 32'h5F5F5F5F;
    'h0757: mem_data <= 32'h2020205F;
    'h0758: mem_data <= 32'h5F5F5F20;
    'h0759: mem_data <= 32'h5F5F5F5F;
    'h075A: mem_data <= 32'h5F5F2020;
    'h075B: mem_data <= 32'h5F5F5F5F;
    'h075C: mem_data <= 32'h5F20205F;
    'h075D: mem_data <= 32'h5F5F5F5F;
    'h075E: mem_data <= 32'h200A5F5F;
    'h075F: mem_data <= 32'h5F5C2020;
    'h0760: mem_data <= 32'h2020205F;
    'h0761: mem_data <= 32'h282F5F5F;
    'h0762: mem_data <= 32'h5F5F2020;
    'h0763: mem_data <= 32'h5C205F5F;
    'h0764: mem_data <= 32'h5F202028;
    'h0765: mem_data <= 32'h205F5F5F;
    'h0766: mem_data <= 32'h2820205C;
    'h0767: mem_data <= 32'h5F5F2020;
    'h0768: mem_data <= 32'h5C205F5F;
    'h0769: mem_data <= 32'h5F202028;
    'h076A: mem_data <= 32'h20205F5F;
    'h076B: mem_data <= 32'h20202829;
    'h076C: mem_data <= 32'h5F5F5F5F;
    'h076D: mem_data <= 32'h200A5C20;
    'h076E: mem_data <= 32'h20202020;
    'h076F: mem_data <= 32'h28202920;
    'h0770: mem_data <= 32'h7C202020;
    'h0771: mem_data <= 32'h20202820;
    'h0772: mem_data <= 32'h2F5C2020;
    'h0773: mem_data <= 32'h2028207C;
    'h0774: mem_data <= 32'h5C202020;
    'h0775: mem_data <= 32'h7C20202F;
    'h0776: mem_data <= 32'h20202820;
    'h0777: mem_data <= 32'h2F5C2020;
    'h0778: mem_data <= 32'h2028207C;
    'h0779: mem_data <= 32'h20292020;
    'h077A: mem_data <= 32'h28207C7C;
    'h077B: mem_data <= 32'h20202020;
    'h077C: mem_data <= 32'h200A2F5C;
    'h077D: mem_data <= 32'h20202020;
    'h077E: mem_data <= 32'h7C207C20;
    'h077F: mem_data <= 32'h7C202020;
    'h0780: mem_data <= 32'h5F5F2820;
    'h0781: mem_data <= 32'h20202020;
    'h0782: mem_data <= 32'h207C207C;
    'h0783: mem_data <= 32'h20202020;
    'h0784: mem_data <= 32'h7C202020;
    'h0785: mem_data <= 32'h5F5F2820;
    'h0786: mem_data <= 32'h205F5F5F;
    'h0787: mem_data <= 32'h207C207C;
    'h0788: mem_data <= 32'h207C2020;
    'h0789: mem_data <= 32'h7C207C7C;
    'h078A: mem_data <= 32'h2020200A;
    'h078B: mem_data <= 32'h7C202020;
    'h078C: mem_data <= 32'h20207C20;
    'h078D: mem_data <= 32'h20207C20;
    'h078E: mem_data <= 32'h20295F5F;
    'h078F: mem_data <= 32'h207C2020;
    'h0790: mem_data <= 32'h5F5F207C;
    'h0791: mem_data <= 32'h20205F5F;
    'h0792: mem_data <= 32'h5F5F2820;
    'h0793: mem_data <= 32'h205F5F5F;
    'h0794: mem_data <= 32'h207C2920;
    'h0795: mem_data <= 32'h2020207C;
    'h0796: mem_data <= 32'h7C7C207C;
    'h0797: mem_data <= 32'h200A7C20;
    'h0798: mem_data <= 32'h20202020;
    'h0799: mem_data <= 32'h7C207C20;
    'h079A: mem_data <= 32'h7C202020;
    'h079B: mem_data <= 32'h20202820;
    'h079C: mem_data <= 32'h20202020;
    'h079D: mem_data <= 32'h207C207C;
    'h079E: mem_data <= 32'h20205F5C;
    'h079F: mem_data <= 32'h20202029;
    'h07A0: mem_data <= 32'h20202020;
    'h07A1: mem_data <= 32'h7C202920;
    'h07A2: mem_data <= 32'h207C207C;
    'h07A3: mem_data <= 32'h207C2020;
    'h07A4: mem_data <= 32'h7C207C7C;
    'h07A5: mem_data <= 32'h2020200A;
    'h07A6: mem_data <= 32'h7C202020;
    'h07A7: mem_data <= 32'h20207C20;
    'h07A8: mem_data <= 32'h29207C20;
    'h07A9: mem_data <= 32'h20202020;
    'h07AA: mem_data <= 32'h207C2020;
    'h07AB: mem_data <= 32'h5F5F5F28;
    'h07AC: mem_data <= 32'h207C2029;
    'h07AD: mem_data <= 32'h5F5C2F20;
    'h07AE: mem_data <= 32'h295F5F5F;
    'h07AF: mem_data <= 32'h207C7C20;
    'h07B0: mem_data <= 32'h5F5F5F28;
    'h07B1: mem_data <= 32'h7C7C2029;
    'h07B2: mem_data <= 32'h5F5F2820;
    'h07B3: mem_data <= 32'h5C2F5F5F;
    'h07B4: mem_data <= 32'h2020200A;
    'h07B5: mem_data <= 32'h29202020;
    'h07B6: mem_data <= 32'h2020285F;
    'h07B7: mem_data <= 32'h202F7C20;
    'h07B8: mem_data <= 32'h20202020;
    'h07B9: mem_data <= 32'h5F282020;
    'h07BA: mem_data <= 32'h5F5F5F5F;
    'h07BB: mem_data <= 32'h20295F5F;
    'h07BC: mem_data <= 32'h5F5F5C20;
    'h07BD: mem_data <= 32'h5F5F5F5F;
    'h07BE: mem_data <= 32'h5F28295F;
    'h07BF: mem_data <= 32'h5F5F5F5F;
    'h07C0: mem_data <= 32'h28295F5F;
    'h07C1: mem_data <= 32'h5F5F5F5F;
    'h07C2: mem_data <= 32'h2F5F5F5F;
    'h07C3: mem_data <= 32'h20410A0A;
    'h07C4: mem_data <= 32'h6B726F66;
    'h07C5: mem_data <= 32'h20666F20;
    'h07C6: mem_data <= 32'h6F636950;
    'h07C7: mem_data <= 32'h20436F53;
    'h07C8: mem_data <= 32'h696C4328;
    'h07C9: mem_data <= 32'h726F6666;
    'h07CA: mem_data <= 32'h6F572064;
    'h07CB: mem_data <= 32'h0A29666C;
    'h07CC: mem_data <= 32'h4F207962;
    'h07CD: mem_data <= 32'h2072616D;
    'h07CE: mem_data <= 32'h656D6F52;
    'h07CF: mem_data <= 32'h000A6172;
    'h07D0: mem_data <= 32'h2020200A;
    'h07D1: mem_data <= 32'h20202020;
    'h07D2: mem_data <= 32'h20202020;
    'h07D3: mem_data <= 32'h20202020;
    'h07D4: mem_data <= 32'h20202020;
    'h07D5: mem_data <= 32'h20202020;
    'h07D6: mem_data <= 32'h20202020;
    'h07D7: mem_data <= 32'h20202020;
    'h07D8: mem_data <= 32'h20202020;
    'h07D9: mem_data <= 32'h20202020;
    'h07DA: mem_data <= 32'h20202020;
    'h07DB: mem_data <= 32'h2D2B2020;
    'h07DC: mem_data <= 32'h202B2D2D;
    'h07DD: mem_data <= 32'h20202020;
    'h07DE: mem_data <= 32'h20202020;
    'h07DF: mem_data <= 32'h20202020;
    'h07E0: mem_data <= 32'h2D2D2D2B;
    'h07E1: mem_data <= 32'h0A2B2D2D;
    'h07E2: mem_data <= 32'h20202020;
    'h07E3: mem_data <= 32'h20202020;
    'h07E4: mem_data <= 32'h20202020;
    'h07E5: mem_data <= 32'h20202020;
    'h07E6: mem_data <= 32'h20202020;
    'h07E7: mem_data <= 32'h20202020;
    'h07E8: mem_data <= 32'h20202020;
    'h07E9: mem_data <= 32'h20202020;
    'h07EA: mem_data <= 32'h20202020;
    'h07EB: mem_data <= 32'h2B202020;
    'h07EC: mem_data <= 32'h2D2D2D2D;
    'h07ED: mem_data <= 32'h57507C2D;
    'h07EE: mem_data <= 32'h2D2D7C52;
    'h07EF: mem_data <= 32'h2D2D2D2D;
    'h07F0: mem_data <= 32'h2D2D2D2D;
    'h07F1: mem_data <= 32'h7C2D2D2D;
    'h07F2: mem_data <= 32'h42535520;
    'h07F3: mem_data <= 32'h2D2D7C20;
    'h07F4: mem_data <= 32'h2B2D2D2D;
    'h07F5: mem_data <= 32'h2020200A;
    'h07F6: mem_data <= 32'h20202020;
    'h07F7: mem_data <= 32'h20202020;
    'h07F8: mem_data <= 32'h20202020;
    'h07F9: mem_data <= 32'h20202020;
    'h07FA: mem_data <= 32'h20202020;
    'h07FB: mem_data <= 32'h20202020;
    'h07FC: mem_data <= 32'h20202020;
    'h07FD: mem_data <= 32'h20202020;
    'h07FE: mem_data <= 32'h20202020;
    'h07FF: mem_data <= 32'h2020207C;
    'h0800: mem_data <= 32'h2D2B2020;
    'h0801: mem_data <= 32'h202B2D2D;
    'h0802: mem_data <= 32'h20202020;
    'h0803: mem_data <= 32'h20202020;
    'h0804: mem_data <= 32'h20202020;
    'h0805: mem_data <= 32'h2D2D2D2B;
    'h0806: mem_data <= 32'h202B2D2D;
    'h0807: mem_data <= 32'h20202020;
    'h0808: mem_data <= 32'h20200A7C;
    'h0809: mem_data <= 32'h20202020;
    'h080A: mem_data <= 32'h20202020;
    'h080B: mem_data <= 32'h20202020;
    'h080C: mem_data <= 32'h20202020;
    'h080D: mem_data <= 32'h20202020;
    'h080E: mem_data <= 32'h20202020;
    'h080F: mem_data <= 32'h20202020;
    'h0810: mem_data <= 32'h20202020;
    'h0811: mem_data <= 32'h20202020;
    'h0812: mem_data <= 32'h20207C20;
    'h0813: mem_data <= 32'h20202020;
    'h0814: mem_data <= 32'h20202020;
    'h0815: mem_data <= 32'h20202020;
    'h0816: mem_data <= 32'h20202020;
    'h0817: mem_data <= 32'h20202020;
    'h0818: mem_data <= 32'h20202020;
    'h0819: mem_data <= 32'h20202020;
    'h081A: mem_data <= 32'h20202020;
    'h081B: mem_data <= 32'h200A7C20;
    'h081C: mem_data <= 32'h20202020;
    'h081D: mem_data <= 32'h20202020;
    'h081E: mem_data <= 32'h20202020;
    'h081F: mem_data <= 32'h4C435320;
    'h0820: mem_data <= 32'h414C535F;
    'h0821: mem_data <= 32'h2F204556;
    'h0822: mem_data <= 32'h4C435320;
    'h0823: mem_data <= 32'h53414D5F;
    'h0824: mem_data <= 32'h20524554;
    'h0825: mem_data <= 32'h207C2020;
    'h0826: mem_data <= 32'h20205858;
    'h0827: mem_data <= 32'h202B2D2B;
    'h0828: mem_data <= 32'h20202020;
    'h0829: mem_data <= 32'h20202020;
    'h082A: mem_data <= 32'h20202020;
    'h082B: mem_data <= 32'h20202020;
    'h082C: mem_data <= 32'h20202020;
    'h082D: mem_data <= 32'hC2202020;
    'h082E: mem_data <= 32'h20B7C2B7;
    'h082F: mem_data <= 32'h20200A7C;
    'h0830: mem_data <= 32'h41445320;
    'h0831: mem_data <= 32'h414C535F;
    'h0832: mem_data <= 32'h2F204556;
    'h0833: mem_data <= 32'h41445320;
    'h0834: mem_data <= 32'h53414D5F;
    'h0835: mem_data <= 32'h20524554;
    'h0836: mem_data <= 32'h5753202F;
    'h0837: mem_data <= 32'h48435449;
    'h0838: mem_data <= 32'h2020335F;
    'h0839: mem_data <= 32'h58207C20;
    'h083A: mem_data <= 32'h7C202058;
    'h083B: mem_data <= 32'h20207C58;
    'h083C: mem_data <= 32'h20202020;
    'h083D: mem_data <= 32'h20202020;
    'h083E: mem_data <= 32'h20202020;
    'h083F: mem_data <= 32'h20202020;
    'h0840: mem_data <= 32'h20202020;
    'h0841: mem_data <= 32'hB7C22020;
    'h0842: mem_data <= 32'h207C2058;
    'h0843: mem_data <= 32'h55532020;
    'h0844: mem_data <= 32'h5F545241;
    'h0845: mem_data <= 32'h200A5854;
    'h0846: mem_data <= 32'h20202020;
    'h0847: mem_data <= 32'h20202020;
    'h0848: mem_data <= 32'h20202020;
    'h0849: mem_data <= 32'h20202020;
    'h084A: mem_data <= 32'h20202020;
    'h084B: mem_data <= 32'h20202020;
    'h084C: mem_data <= 32'h53202020;
    'h084D: mem_data <= 32'h43544957;
    'h084E: mem_data <= 32'h20325F48;
    'h084F: mem_data <= 32'h207C2020;
    'h0850: mem_data <= 32'hB7C2B7C2;
    'h0851: mem_data <= 32'h587C2020;
    'h0852: mem_data <= 32'h2020207C;
    'h0853: mem_data <= 32'h20202020;
    'h0854: mem_data <= 32'h20202020;
    'h0855: mem_data <= 32'h4C202020;
    'h0856: mem_data <= 32'h20374445;
    'h0857: mem_data <= 32'h207D587B;
    'h0858: mem_data <= 32'h58B7C220;
    'h0859: mem_data <= 32'h20207C20;
    'h085A: mem_data <= 32'h44454C20;
    'h085B: mem_data <= 32'h2F20375F;
    'h085C: mem_data <= 32'h41555320;
    'h085D: mem_data <= 32'h525F5452;
    'h085E: mem_data <= 32'h20200A58;
    'h085F: mem_data <= 32'h20202020;
    'h0860: mem_data <= 32'h20202020;
    'h0861: mem_data <= 32'h20202020;
    'h0862: mem_data <= 32'h20202020;
    'h0863: mem_data <= 32'h20202020;
    'h0864: mem_data <= 32'h20202020;
    'h0865: mem_data <= 32'h57532020;
    'h0866: mem_data <= 32'h48435449;
    'h0867: mem_data <= 32'h2020315F;
    'h0868: mem_data <= 32'hC2207C20;
    'h0869: mem_data <= 32'h20B7C2B7;
    'h086A: mem_data <= 32'h7C587C20;
    'h086B: mem_data <= 32'h20202020;
    'h086C: mem_data <= 32'h20202020;
    'h086D: mem_data <= 32'h20202020;
    'h086E: mem_data <= 32'h454C2020;
    'h086F: mem_data <= 32'h7B203644;
    'h0870: mem_data <= 32'h20207D58;
    'h0871: mem_data <= 32'hB7C2B7C2;
    'h0872: mem_data <= 32'h20207C20;
    'h0873: mem_data <= 32'h44454C20;
    'h0874: mem_data <= 32'h200A365F;
    'h0875: mem_data <= 32'h20202020;
    'h0876: mem_data <= 32'h20202020;
    'h0877: mem_data <= 32'h20202020;
    'h0878: mem_data <= 32'h20202020;
    'h0879: mem_data <= 32'h20202020;
    'h087A: mem_data <= 32'h20202020;
    'h087B: mem_data <= 32'h53202020;
    'h087C: mem_data <= 32'h43544957;
    'h087D: mem_data <= 32'h20305F48;
    'h087E: mem_data <= 32'h207C2020;
    'h087F: mem_data <= 32'hB7C2B7C2;
    'h0880: mem_data <= 32'h587C2020;
    'h0881: mem_data <= 32'h2020207C;
    'h0882: mem_data <= 32'h20202020;
    'h0883: mem_data <= 32'h20202020;
    'h0884: mem_data <= 32'h4C202020;
    'h0885: mem_data <= 32'h20354445;
    'h0886: mem_data <= 32'h207D587B;
    'h0887: mem_data <= 32'hC2B7C220;
    'h0888: mem_data <= 32'h207C20B7;
    'h0889: mem_data <= 32'h454C2020;
    'h088A: mem_data <= 32'h0A355F44;
    'h088B: mem_data <= 32'h20202020;
    'h088C: mem_data <= 32'h20202020;
    'h088D: mem_data <= 32'h20202020;
    'h088E: mem_data <= 32'h20202020;
    'h088F: mem_data <= 32'h20202020;
    'h0890: mem_data <= 32'h20202020;
    'h0891: mem_data <= 32'h20202020;
    'h0892: mem_data <= 32'h63562020;
    'h0893: mem_data <= 32'h33703363;
    'h0894: mem_data <= 32'h7C202020;
    'h0895: mem_data <= 32'h58B7C220;
    'h0896: mem_data <= 32'h2D2B2020;
    'h0897: mem_data <= 32'h2020202B;
    'h0898: mem_data <= 32'h20202020;
    'h0899: mem_data <= 32'h20202020;
    'h089A: mem_data <= 32'h4C202020;
    'h089B: mem_data <= 32'h20344445;
    'h089C: mem_data <= 32'h207D587B;
    'h089D: mem_data <= 32'h20585820;
    'h089E: mem_data <= 32'h2020207C;
    'h089F: mem_data <= 32'h5F44454C;
    'h08A0: mem_data <= 32'h202F2034;
    'h08A1: mem_data <= 32'h35636356;
    'h08A2: mem_data <= 32'h47202F20;
    'h08A3: mem_data <= 32'h200A444E;
    'h08A4: mem_data <= 32'h20202020;
    'h08A5: mem_data <= 32'h20202020;
    'h08A6: mem_data <= 32'h20202020;
    'h08A7: mem_data <= 32'h20202020;
    'h08A8: mem_data <= 32'h20202020;
    'h08A9: mem_data <= 32'h20202020;
    'h08AA: mem_data <= 32'h20202020;
    'h08AB: mem_data <= 32'h20202020;
    'h08AC: mem_data <= 32'h20202020;
    'h08AD: mem_data <= 32'h207C2020;
    'h08AE: mem_data <= 32'hB7C2B7C2;
    'h08AF: mem_data <= 32'h20202020;
    'h08B0: mem_data <= 32'h20202020;
    'h08B1: mem_data <= 32'h20202020;
    'h08B2: mem_data <= 32'h20202020;
    'h08B3: mem_data <= 32'h4C202020;
    'h08B4: mem_data <= 32'h20334445;
    'h08B5: mem_data <= 32'h207D587B;
    'h08B6: mem_data <= 32'hC2B7C220;
    'h08B7: mem_data <= 32'h207C20B7;
    'h08B8: mem_data <= 32'h454C2020;
    'h08B9: mem_data <= 32'h0A335F44;
    'h08BA: mem_data <= 32'h20202020;
    'h08BB: mem_data <= 32'h20202020;
    'h08BC: mem_data <= 32'h20202020;
    'h08BD: mem_data <= 32'h20202020;
    'h08BE: mem_data <= 32'h20202020;
    'h08BF: mem_data <= 32'h20202020;
    'h08C0: mem_data <= 32'h20202020;
    'h08C1: mem_data <= 32'h20202020;
    'h08C2: mem_data <= 32'h20202020;
    'h08C3: mem_data <= 32'h7C202020;
    'h08C4: mem_data <= 32'hC2B7C220;
    'h08C5: mem_data <= 32'h202020B7;
    'h08C6: mem_data <= 32'h20202020;
    'h08C7: mem_data <= 32'h20202020;
    'h08C8: mem_data <= 32'h20202020;
    'h08C9: mem_data <= 32'h20202020;
    'h08CA: mem_data <= 32'h3244454C;
    'h08CB: mem_data <= 32'h7D587B20;
    'h08CC: mem_data <= 32'hB7C22020;
    'h08CD: mem_data <= 32'h7C20B7C2;
    'h08CE: mem_data <= 32'h4C202020;
    'h08CF: mem_data <= 32'h325F4445;
    'h08D0: mem_data <= 32'h2020200A;
    'h08D1: mem_data <= 32'h20202020;
    'h08D2: mem_data <= 32'h20202020;
    'h08D3: mem_data <= 32'h20202020;
    'h08D4: mem_data <= 32'h20202020;
    'h08D5: mem_data <= 32'h20202020;
    'h08D6: mem_data <= 32'h20202020;
    'h08D7: mem_data <= 32'h20202020;
    'h08D8: mem_data <= 32'h20202020;
    'h08D9: mem_data <= 32'h20202020;
    'h08DA: mem_data <= 32'hB7C2207C;
    'h08DB: mem_data <= 32'h2020B7C2;
    'h08DC: mem_data <= 32'h20202020;
    'h08DD: mem_data <= 32'h20202020;
    'h08DE: mem_data <= 32'h20202020;
    'h08DF: mem_data <= 32'h20202020;
    'h08E0: mem_data <= 32'h44454C20;
    'h08E1: mem_data <= 32'h587B2031;
    'h08E2: mem_data <= 32'hC220207D;
    'h08E3: mem_data <= 32'h20B7C2B7;
    'h08E4: mem_data <= 32'h2020207C;
    'h08E5: mem_data <= 32'h5F44454C;
    'h08E6: mem_data <= 32'h20200A31;
    'h08E7: mem_data <= 32'h20202020;
    'h08E8: mem_data <= 32'h20202020;
    'h08E9: mem_data <= 32'h20202020;
    'h08EA: mem_data <= 32'h20202020;
    'h08EB: mem_data <= 32'h20202020;
    'h08EC: mem_data <= 32'h20202020;
    'h08ED: mem_data <= 32'h20202020;
    'h08EE: mem_data <= 32'h20202020;
    'h08EF: mem_data <= 32'h20202020;
    'h08F0: mem_data <= 32'hC2207C20;
    'h08F1: mem_data <= 32'h20B7C2B7;
    'h08F2: mem_data <= 32'h20202020;
    'h08F3: mem_data <= 32'h20202020;
    'h08F4: mem_data <= 32'h20202020;
    'h08F5: mem_data <= 32'h20202020;
    'h08F6: mem_data <= 32'h454C2020;
    'h08F7: mem_data <= 32'h7B203044;
    'h08F8: mem_data <= 32'h20207D58;
    'h08F9: mem_data <= 32'hB7C2B7C2;
    'h08FA: mem_data <= 32'h20207C20;
    'h08FB: mem_data <= 32'h44454C20;
    'h08FC: mem_data <= 32'h200A305F;
    'h08FD: mem_data <= 32'h20202020;
    'h08FE: mem_data <= 32'h20202020;
    'h08FF: mem_data <= 32'h20202020;
    'h0900: mem_data <= 32'h20202020;
    'h0901: mem_data <= 32'h20202020;
    'h0902: mem_data <= 32'h20202020;
    'h0903: mem_data <= 32'h20202020;
    'h0904: mem_data <= 32'h20202020;
    'h0905: mem_data <= 32'h20202020;
    'h0906: mem_data <= 32'h207C2020;
    'h0907: mem_data <= 32'hB7C2B7C2;
    'h0908: mem_data <= 32'h20202020;
    'h0909: mem_data <= 32'h20202020;
    'h090A: mem_data <= 32'h20202020;
    'h090B: mem_data <= 32'h20202020;
    'h090C: mem_data <= 32'h20202020;
    'h090D: mem_data <= 32'h20202020;
    'h090E: mem_data <= 32'h20202020;
    'h090F: mem_data <= 32'hC2B7C220;
    'h0910: mem_data <= 32'h0A7C20B7;
    'h0911: mem_data <= 32'h20202020;
    'h0912: mem_data <= 32'h20202020;
    'h0913: mem_data <= 32'h20202020;
    'h0914: mem_data <= 32'h20202020;
    'h0915: mem_data <= 32'h20202020;
    'h0916: mem_data <= 32'h20202020;
    'h0917: mem_data <= 32'h20202020;
    'h0918: mem_data <= 32'h20202020;
    'h0919: mem_data <= 32'h20202020;
    'h091A: mem_data <= 32'h7C202020;
    'h091B: mem_data <= 32'hC2B7C220;
    'h091C: mem_data <= 32'h202020B7;
    'h091D: mem_data <= 32'h2D2D2B20;
    'h091E: mem_data <= 32'h2D2D2D2D;
    'h091F: mem_data <= 32'h2D2D2D2D;
    'h0920: mem_data <= 32'h2D2D2D2D;
    'h0921: mem_data <= 32'h20202B2D;
    'h0922: mem_data <= 32'h20202020;
    'h0923: mem_data <= 32'hB7C22020;
    'h0924: mem_data <= 32'h7C20B7C2;
    'h0925: mem_data <= 32'h2020200A;
    'h0926: mem_data <= 32'h20202020;
    'h0927: mem_data <= 32'h20202020;
    'h0928: mem_data <= 32'h20202020;
    'h0929: mem_data <= 32'h20202020;
    'h092A: mem_data <= 32'h20202020;
    'h092B: mem_data <= 32'h20202020;
    'h092C: mem_data <= 32'h20202020;
    'h092D: mem_data <= 32'h20202020;
    'h092E: mem_data <= 32'h20202020;
    'h092F: mem_data <= 32'hB7C2207C;
    'h0930: mem_data <= 32'h2020B7C2;
    'h0931: mem_data <= 32'h207C2020;
    'h0932: mem_data <= 32'h20202020;
    'h0933: mem_data <= 32'h20202020;
    'h0934: mem_data <= 32'h20202020;
    'h0935: mem_data <= 32'h207C2020;
    'h0936: mem_data <= 32'h20202020;
    'h0937: mem_data <= 32'hC2202020;
    'h0938: mem_data <= 32'h20B7C2B7;
    'h0939: mem_data <= 32'h20200A7C;
    'h093A: mem_data <= 32'h20202020;
    'h093B: mem_data <= 32'h20202020;
    'h093C: mem_data <= 32'h20202020;
    'h093D: mem_data <= 32'h20202020;
    'h093E: mem_data <= 32'h20202020;
    'h093F: mem_data <= 32'h20202020;
    'h0940: mem_data <= 32'h20202020;
    'h0941: mem_data <= 32'h20202020;
    'h0942: mem_data <= 32'h20202020;
    'h0943: mem_data <= 32'hC2207C20;
    'h0944: mem_data <= 32'h20B7C2B7;
    'h0945: mem_data <= 32'h7C202020;
    'h0946: mem_data <= 32'h20202020;
    'h0947: mem_data <= 32'h20202020;
    'h0948: mem_data <= 32'h20202020;
    'h0949: mem_data <= 32'h7C202020;
    'h094A: mem_data <= 32'h2B202020;
    'h094B: mem_data <= 32'h20202B2D;
    'h094C: mem_data <= 32'hB7C2B7C2;
    'h094D: mem_data <= 32'h200A7C20;
    'h094E: mem_data <= 32'h20202020;
    'h094F: mem_data <= 32'h20202020;
    'h0950: mem_data <= 32'h20202020;
    'h0951: mem_data <= 32'h20202020;
    'h0952: mem_data <= 32'h20202020;
    'h0953: mem_data <= 32'h20202020;
    'h0954: mem_data <= 32'h20202020;
    'h0955: mem_data <= 32'h20202020;
    'h0956: mem_data <= 32'h20202020;
    'h0957: mem_data <= 32'h207C2020;
    'h0958: mem_data <= 32'hB7C2B7C2;
    'h0959: mem_data <= 32'h20202020;
    'h095A: mem_data <= 32'h4320207C;
    'h095B: mem_data <= 32'h6F6C6379;
    'h095C: mem_data <= 32'h2020656E;
    'h095D: mem_data <= 32'h20205649;
    'h095E: mem_data <= 32'h2020207C;
    'h095F: mem_data <= 32'h207C587C;
    'h0960: mem_data <= 32'hB7C25820;
    'h0961: mem_data <= 32'h20207C20;
    'h0962: mem_data <= 32'h54554220;
    'h0963: mem_data <= 32'h5F4E4F54;
    'h0964: mem_data <= 32'h202F2031;
    'h0965: mem_data <= 32'h33636356;
    'h0966: mem_data <= 32'h200A3370;
    'h0967: mem_data <= 32'h20202020;
    'h0968: mem_data <= 32'h20202020;
    'h0969: mem_data <= 32'h20202020;
    'h096A: mem_data <= 32'h20202020;
    'h096B: mem_data <= 32'h20202020;
    'h096C: mem_data <= 32'h20202020;
    'h096D: mem_data <= 32'h20202020;
    'h096E: mem_data <= 32'h20202020;
    'h096F: mem_data <= 32'h20202020;
    'h0970: mem_data <= 32'h207C2020;
    'h0971: mem_data <= 32'hB7C2B7C2;
    'h0972: mem_data <= 32'h20202020;
    'h0973: mem_data <= 32'h2020207C;
    'h0974: mem_data <= 32'h20202020;
    'h0975: mem_data <= 32'h20202020;
    'h0976: mem_data <= 32'h20202020;
    'h0977: mem_data <= 32'h2020207C;
    'h0978: mem_data <= 32'h202B2D2B;
    'h0979: mem_data <= 32'hC2B7C220;
    'h097A: mem_data <= 32'h0A7C20B7;
    'h097B: mem_data <= 32'h20202020;
    'h097C: mem_data <= 32'h20202020;
    'h097D: mem_data <= 32'h20202020;
    'h097E: mem_data <= 32'h20202020;
    'h097F: mem_data <= 32'h20202020;
    'h0980: mem_data <= 32'h20202020;
    'h0981: mem_data <= 32'h20202020;
    'h0982: mem_data <= 32'h20202020;
    'h0983: mem_data <= 32'h20202020;
    'h0984: mem_data <= 32'h7C202020;
    'h0985: mem_data <= 32'hC2B7C220;
    'h0986: mem_data <= 32'h202020B7;
    'h0987: mem_data <= 32'h45207C20;
    'h0988: mem_data <= 32'h45433450;
    'h0989: mem_data <= 32'h31463232;
    'h098A: mem_data <= 32'h4E364337;
    'h098B: mem_data <= 32'h20207C20;
    'h098C: mem_data <= 32'h20202020;
    'h098D: mem_data <= 32'hB7C22020;
    'h098E: mem_data <= 32'h7C20B7C2;
    'h098F: mem_data <= 32'h2020200A;
    'h0990: mem_data <= 32'h20202020;
    'h0991: mem_data <= 32'h20202020;
    'h0992: mem_data <= 32'h20202020;
    'h0993: mem_data <= 32'h20202020;
    'h0994: mem_data <= 32'h20202020;
    'h0995: mem_data <= 32'h20202020;
    'h0996: mem_data <= 32'h20202020;
    'h0997: mem_data <= 32'h20202020;
    'h0998: mem_data <= 32'h20202020;
    'h0999: mem_data <= 32'hB7C2207C;
    'h099A: mem_data <= 32'h2020B7C2;
    'h099B: mem_data <= 32'h207C2020;
    'h099C: mem_data <= 32'h20202020;
    'h099D: mem_data <= 32'h20202020;
    'h099E: mem_data <= 32'h20202020;
    'h099F: mem_data <= 32'h207C2020;
    'h09A0: mem_data <= 32'h2D2B2020;
    'h09A1: mem_data <= 32'hC220202B;
    'h09A2: mem_data <= 32'h20B7C2B7;
    'h09A3: mem_data <= 32'h20200A7C;
    'h09A4: mem_data <= 32'h20202020;
    'h09A5: mem_data <= 32'h20202020;
    'h09A6: mem_data <= 32'h20202020;
    'h09A7: mem_data <= 32'h20202020;
    'h09A8: mem_data <= 32'h20202020;
    'h09A9: mem_data <= 32'h20202020;
    'h09AA: mem_data <= 32'h20202020;
    'h09AB: mem_data <= 32'h20202020;
    'h09AC: mem_data <= 32'h20202020;
    'h09AD: mem_data <= 32'hC2207C20;
    'h09AE: mem_data <= 32'h20B7C2B7;
    'h09AF: mem_data <= 32'h7C202020;
    'h09B0: mem_data <= 32'h20202020;
    'h09B1: mem_data <= 32'h20202020;
    'h09B2: mem_data <= 32'h20202020;
    'h09B3: mem_data <= 32'h7C202020;
    'h09B4: mem_data <= 32'h7C202020;
    'h09B5: mem_data <= 32'h20207C58;
    'h09B6: mem_data <= 32'hB7C2B7C2;
    'h09B7: mem_data <= 32'h20207C20;
    'h09B8: mem_data <= 32'h54554220;
    'h09B9: mem_data <= 32'h5F4E4F54;
    'h09BA: mem_data <= 32'h20200A30;
    'h09BB: mem_data <= 32'h20202020;
    'h09BC: mem_data <= 32'h20202020;
    'h09BD: mem_data <= 32'h20202020;
    'h09BE: mem_data <= 32'h20202020;
    'h09BF: mem_data <= 32'h20202020;
    'h09C0: mem_data <= 32'h20202020;
    'h09C1: mem_data <= 32'h20202020;
    'h09C2: mem_data <= 32'h20202020;
    'h09C3: mem_data <= 32'h20202020;
    'h09C4: mem_data <= 32'hC2207C20;
    'h09C5: mem_data <= 32'h20B7C2B7;
    'h09C6: mem_data <= 32'h2B202020;
    'h09C7: mem_data <= 32'h2D2D2D2D;
    'h09C8: mem_data <= 32'h2D2D2D2D;
    'h09C9: mem_data <= 32'h2D2D2D2D;
    'h09CA: mem_data <= 32'h2B2D2D2D;
    'h09CB: mem_data <= 32'h2B202020;
    'h09CC: mem_data <= 32'h20202B2D;
    'h09CD: mem_data <= 32'hB7C2B7C2;
    'h09CE: mem_data <= 32'h200A7C20;
    'h09CF: mem_data <= 32'h20202020;
    'h09D0: mem_data <= 32'h20202020;
    'h09D1: mem_data <= 32'h20202020;
    'h09D2: mem_data <= 32'h20202020;
    'h09D3: mem_data <= 32'h20202020;
    'h09D4: mem_data <= 32'h20202020;
    'h09D5: mem_data <= 32'h20202020;
    'h09D6: mem_data <= 32'h20202020;
    'h09D7: mem_data <= 32'h20202020;
    'h09D8: mem_data <= 32'h207C2020;
    'h09D9: mem_data <= 32'h20202020;
    'h09DA: mem_data <= 32'h20202020;
    'h09DB: mem_data <= 32'h20202020;
    'h09DC: mem_data <= 32'h20202020;
    'h09DD: mem_data <= 32'h20202020;
    'h09DE: mem_data <= 32'h20202020;
    'h09DF: mem_data <= 32'h20202020;
    'h09E0: mem_data <= 32'h20202020;
    'h09E1: mem_data <= 32'h0A7C2020;
    'h09E2: mem_data <= 32'h20202020;
    'h09E3: mem_data <= 32'h20202020;
    'h09E4: mem_data <= 32'h20202020;
    'h09E5: mem_data <= 32'h20202020;
    'h09E6: mem_data <= 32'h20202020;
    'h09E7: mem_data <= 32'h20202020;
    'h09E8: mem_data <= 32'h20202020;
    'h09E9: mem_data <= 32'h20202020;
    'h09EA: mem_data <= 32'h20202020;
    'h09EB: mem_data <= 32'h7C202020;
    'h09EC: mem_data <= 32'h20202020;
    'h09ED: mem_data <= 32'h20B7C220;
    'h09EE: mem_data <= 32'hC220B7C2;
    'h09EF: mem_data <= 32'hB7C220B7;
    'h09F0: mem_data <= 32'h20B7C220;
    'h09F1: mem_data <= 32'hC220B7C2;
    'h09F2: mem_data <= 32'hB7C220B7;
    'h09F3: mem_data <= 32'h20B7C220;
    'h09F4: mem_data <= 32'hC220B7C2;
    'h09F5: mem_data <= 32'hB7C220B7;
    'h09F6: mem_data <= 32'h20B7C220;
    'h09F7: mem_data <= 32'h20202020;
    'h09F8: mem_data <= 32'h20200A7C;
    'h09F9: mem_data <= 32'h20202020;
    'h09FA: mem_data <= 32'h20202020;
    'h09FB: mem_data <= 32'h20202020;
    'h09FC: mem_data <= 32'h20202020;
    'h09FD: mem_data <= 32'h20202020;
    'h09FE: mem_data <= 32'h20202020;
    'h09FF: mem_data <= 32'h20202020;
    'h0A00: mem_data <= 32'h20202020;
    'h0A01: mem_data <= 32'h20202020;
    'h0A02: mem_data <= 32'h20207C20;
    'h0A03: mem_data <= 32'hC2202020;
    'h0A04: mem_data <= 32'hB7C220B7;
    'h0A05: mem_data <= 32'h20B7C220;
    'h0A06: mem_data <= 32'hC220B7C2;
    'h0A07: mem_data <= 32'hB7C220B7;
    'h0A08: mem_data <= 32'h20B7C220;
    'h0A09: mem_data <= 32'hC220B7C2;
    'h0A0A: mem_data <= 32'hB7C220B7;
    'h0A0B: mem_data <= 32'h20B7C220;
    'h0A0C: mem_data <= 32'hC220B7C2;
    'h0A0D: mem_data <= 32'h202020B7;
    'h0A0E: mem_data <= 32'h0A7C2020;
    'h0A0F: mem_data <= 32'h20202020;
    'h0A10: mem_data <= 32'h20202020;
    'h0A11: mem_data <= 32'h20202020;
    'h0A12: mem_data <= 32'h20202020;
    'h0A13: mem_data <= 32'h20202020;
    'h0A14: mem_data <= 32'h20202020;
    'h0A15: mem_data <= 32'h20202020;
    'h0A16: mem_data <= 32'h20202020;
    'h0A17: mem_data <= 32'h20202020;
    'h0A18: mem_data <= 32'h2B202020;
    'h0A19: mem_data <= 32'h2D2D2D2D;
    'h0A1A: mem_data <= 32'h2D2D2D2D;
    'h0A1B: mem_data <= 32'h2D2D2D2D;
    'h0A1C: mem_data <= 32'h2D2D2D2D;
    'h0A1D: mem_data <= 32'h2D2D2D2D;
    'h0A1E: mem_data <= 32'h2D2D2D2D;
    'h0A1F: mem_data <= 32'h2D2D2D2D;
    'h0A20: mem_data <= 32'h2D2D2D2D;
    'h0A21: mem_data <= 32'h2B2D2D2D;
    'h0A22: mem_data <= 32'h00000A0A;
    'h0A23: mem_data <= 32'h204E4950;
    'h0A24: mem_data <= 32'h7473694C;
    'h0A25: mem_data <= 32'h200A0A3A;
    'h0A26: mem_data <= 32'h32492020;
    'h0A27: mem_data <= 32'h20200A43;
    'h0A28: mem_data <= 32'h20202020;
    'h0A29: mem_data <= 32'h2034314A;
    'h0A2A: mem_data <= 32'h2D202020;
    'h0A2B: mem_data <= 32'h4C435320;
    'h0A2C: mem_data <= 32'h414C535F;
    'h0A2D: mem_data <= 32'h200A4556;
    'h0A2E: mem_data <= 32'h20202020;
    'h0A2F: mem_data <= 32'h33314A20;
    'h0A30: mem_data <= 32'h20202020;
    'h0A31: mem_data <= 32'h4353202D;
    'h0A32: mem_data <= 32'h414D5F4C;
    'h0A33: mem_data <= 32'h52455453;
    'h0A34: mem_data <= 32'h2020200A;
    'h0A35: mem_data <= 32'h4B202020;
    'h0A36: mem_data <= 32'h20203531;
    'h0A37: mem_data <= 32'h202D2020;
    'h0A38: mem_data <= 32'h5F414453;
    'h0A39: mem_data <= 32'h56414C53;
    'h0A3A: mem_data <= 32'h20200A45;
    'h0A3B: mem_data <= 32'h20202020;
    'h0A3C: mem_data <= 32'h2036314A;
    'h0A3D: mem_data <= 32'h2D202020;
    'h0A3E: mem_data <= 32'h41445320;
    'h0A3F: mem_data <= 32'h53414D5F;
    'h0A40: mem_data <= 32'h0A524554;
    'h0A41: mem_data <= 32'h20202020;
    'h0A42: mem_data <= 32'h63562020;
    'h0A43: mem_data <= 32'h33703363;
    'h0A44: mem_data <= 32'h50202D20;
    'h0A45: mem_data <= 32'h204C4C55;
    'h0A46: mem_data <= 32'h52205055;
    'h0A47: mem_data <= 32'h53495345;
    'h0A48: mem_data <= 32'h20524F54;
    'h0A49: mem_data <= 32'h0A0A4B31;
    'h0A4A: mem_data <= 32'h53202020;
    'h0A4B: mem_data <= 32'h555F5359;
    'h0A4C: mem_data <= 32'h0A545241;
    'h0A4D: mem_data <= 32'h20202020;
    'h0A4E: mem_data <= 32'h33412020;
    'h0A4F: mem_data <= 32'h20202020;
    'h0A50: mem_data <= 32'h53202D20;
    'h0A51: mem_data <= 32'h54524155;
    'h0A52: mem_data <= 32'h0A58525F;
    'h0A53: mem_data <= 32'h20202020;
    'h0A54: mem_data <= 32'h33432020;
    'h0A55: mem_data <= 32'h20202020;
    'h0A56: mem_data <= 32'h53202D20;
    'h0A57: mem_data <= 32'h54524155;
    'h0A58: mem_data <= 32'h0A58545F;
    'h0A59: mem_data <= 32'h2020200A;
    'h0A5A: mem_data <= 32'h5344454C;
    'h0A5B: mem_data <= 32'h2020200A;
    'h0A5C: mem_data <= 32'h41202020;
    'h0A5D: mem_data <= 32'h20203531;
    'h0A5E: mem_data <= 32'h202D2020;
    'h0A5F: mem_data <= 32'h5F44454C;
    'h0A60: mem_data <= 32'h20200A30;
    'h0A61: mem_data <= 32'h20202020;
    'h0A62: mem_data <= 32'h20333141;
    'h0A63: mem_data <= 32'h2D202020;
    'h0A64: mem_data <= 32'h44454C20;
    'h0A65: mem_data <= 32'h200A315F;
    'h0A66: mem_data <= 32'h20202020;
    'h0A67: mem_data <= 32'h33314220;
    'h0A68: mem_data <= 32'h20202020;
    'h0A69: mem_data <= 32'h454C202D;
    'h0A6A: mem_data <= 32'h0A325F44;
    'h0A6B: mem_data <= 32'h20202020;
    'h0A6C: mem_data <= 32'h31412020;
    'h0A6D: mem_data <= 32'h20202031;
    'h0A6E: mem_data <= 32'h4C202D20;
    'h0A6F: mem_data <= 32'h335F4445;
    'h0A70: mem_data <= 32'h2020200A;
    'h0A71: mem_data <= 32'h44202020;
    'h0A72: mem_data <= 32'h20202031;
    'h0A73: mem_data <= 32'h202D2020;
    'h0A74: mem_data <= 32'h5F44454C;
    'h0A75: mem_data <= 32'h20200A34;
    'h0A76: mem_data <= 32'h20202020;
    'h0A77: mem_data <= 32'h20203346;
    'h0A78: mem_data <= 32'h2D202020;
    'h0A79: mem_data <= 32'h44454C20;
    'h0A7A: mem_data <= 32'h200A355F;
    'h0A7B: mem_data <= 32'h20202020;
    'h0A7C: mem_data <= 32'h20314220;
    'h0A7D: mem_data <= 32'h20202020;
    'h0A7E: mem_data <= 32'h454C202D;
    'h0A7F: mem_data <= 32'h0A365F44;
    'h0A80: mem_data <= 32'h20202020;
    'h0A81: mem_data <= 32'h334C2020;
    'h0A82: mem_data <= 32'h20202020;
    'h0A83: mem_data <= 32'h4C202D20;
    'h0A84: mem_data <= 32'h375F4445;
    'h0A85: mem_data <= 32'h20200A0A;
    'h0A86: mem_data <= 32'h54554220;
    'h0A87: mem_data <= 32'h534E4F54;
    'h0A88: mem_data <= 32'h2020200A;
    'h0A89: mem_data <= 32'h4A202020;
    'h0A8A: mem_data <= 32'h20203531;
    'h0A8B: mem_data <= 32'h202D2020;
    'h0A8C: mem_data <= 32'h54545542;
    'h0A8D: mem_data <= 32'h305F4E4F;
    'h0A8E: mem_data <= 32'h2020200A;
    'h0A8F: mem_data <= 32'h45202020;
    'h0A90: mem_data <= 32'h20202031;
    'h0A91: mem_data <= 32'h202D2020;
    'h0A92: mem_data <= 32'h54545542;
    'h0A93: mem_data <= 32'h315F4E4F;
    'h0A94: mem_data <= 32'h20200A0A;
    'h0A95: mem_data <= 32'h49575320;
    'h0A96: mem_data <= 32'h45484354;
    'h0A97: mem_data <= 32'h20200A53;
    'h0A98: mem_data <= 32'h20202020;
    'h0A99: mem_data <= 32'h2020314D;
    'h0A9A: mem_data <= 32'h2D202020;
    'h0A9B: mem_data <= 32'h49575320;
    'h0A9C: mem_data <= 32'h5F484354;
    'h0A9D: mem_data <= 32'h20200A30;
    'h0A9E: mem_data <= 32'h20202020;
    'h0A9F: mem_data <= 32'h20203854;
    'h0AA0: mem_data <= 32'h2D202020;
    'h0AA1: mem_data <= 32'h49575320;
    'h0AA2: mem_data <= 32'h5F484354;
    'h0AA3: mem_data <= 32'h20200A31;
    'h0AA4: mem_data <= 32'h20202020;
    'h0AA5: mem_data <= 32'h20203942;
    'h0AA6: mem_data <= 32'h2D202020;
    'h0AA7: mem_data <= 32'h49575320;
    'h0AA8: mem_data <= 32'h5F484354;
    'h0AA9: mem_data <= 32'h20200A32;
    'h0AAA: mem_data <= 32'h20202020;
    'h0AAB: mem_data <= 32'h2035314D;
    'h0AAC: mem_data <= 32'h2D202020;
    'h0AAD: mem_data <= 32'h49575320;
    'h0AAE: mem_data <= 32'h5F484354;
    'h0AAF: mem_data <= 32'h000A0A33;
    'h0AB0: mem_data <= 32'h20200A0A;
    'h0AB1: mem_data <= 32'h5D315B20;
    'h0AB2: mem_data <= 32'h6E695020;
    'h0AB3: mem_data <= 32'h2074756F;
    'h0AB4: mem_data <= 32'h0A70614D;
    'h0AB5: mem_data <= 32'h5B202020;
    'h0AB6: mem_data <= 32'h50205D32;
    'h0AB7: mem_data <= 32'h756F6E69;
    'h0AB8: mem_data <= 32'h694C2074;
    'h0AB9: mem_data <= 32'h200A7473;
    'h0ABA: mem_data <= 32'h335B2020;
    'h0ABB: mem_data <= 32'h5047205D;
    'h0ABC: mem_data <= 32'h74204F49;
    'h0ABD: mem_data <= 32'h62747365;
    'h0ABE: mem_data <= 32'h68636E65;
    'h0ABF: mem_data <= 32'h2020200A;
    'h0AC0: mem_data <= 32'h205D345B;
    'h0AC1: mem_data <= 32'h20433249;
    'h0AC2: mem_data <= 32'h74736574;
    'h0AC3: mem_data <= 32'h636E6562;
    'h0AC4: mem_data <= 32'h20200A68;
    'h0AC5: mem_data <= 32'h5D355B20;
    'h0AC6: mem_data <= 32'h49505320;
    'h0AC7: mem_data <= 32'h73657420;
    'h0AC8: mem_data <= 32'h6E656274;
    'h0AC9: mem_data <= 32'h0A0A6863;
    'h0ACA: mem_data <= 32'h00000000;
    'h0ACB: mem_data <= 32'h656C6553;
    'h0ACC: mem_data <= 32'h6F207463;
    'h0ACD: mem_data <= 32'h6F697470;
    'h0ACE: mem_data <= 32'h00203E6E;
    'h0ACF: mem_data <= 32'h0010153C;
    'h0AD0: mem_data <= 32'h0010154C;
    'h0AD1: mem_data <= 32'h0010155C;
    'h0AD2: mem_data <= 32'h00101568;
    'h0AD3: mem_data <= 32'h00101574;
    'h0AD4: mem_data <= 32'h20200A0A;
    'h0AD5: mem_data <= 32'h5D315B20;
    'h0AD6: mem_data <= 32'h6E755220;
    'h0AD7: mem_data <= 32'h44454C20;
    'h0AD8: mem_data <= 32'h73657420;
    'h0AD9: mem_data <= 32'h6E656274;
    'h0ADA: mem_data <= 32'h200A6863;
    'h0ADB: mem_data <= 32'h325B2020;
    'h0ADC: mem_data <= 32'h7552205D;
    'h0ADD: mem_data <= 32'h5542206E;
    'h0ADE: mem_data <= 32'h4E4F5454;
    'h0ADF: mem_data <= 32'h6E612053;
    'h0AE0: mem_data <= 32'h57532064;
    'h0AE1: mem_data <= 32'h48435449;
    'h0AE2: mem_data <= 32'h74205345;
    'h0AE3: mem_data <= 32'h62747365;
    'h0AE4: mem_data <= 32'h68636E65;
    'h0AE5: mem_data <= 32'h2020200A;
    'h0AE6: mem_data <= 32'h205D725B;
    'h0AE7: mem_data <= 32'h75746552;
    'h0AE8: mem_data <= 32'h74206E72;
    'h0AE9: mem_data <= 32'h616D206F;
    'h0AEA: mem_data <= 32'h6D206E69;
    'h0AEB: mem_data <= 32'h0A756E65;
    'h0AEC: mem_data <= 32'h0000000A;
    'h0AED: mem_data <= 32'h656C6553;
    'h0AEE: mem_data <= 32'h6D207463;
    'h0AEF: mem_data <= 32'h3E65646F;
    'h0AF0: mem_data <= 32'h00000020;
    'h0AF1: mem_data <= 32'h20200A0A;
    'h0AF2: mem_data <= 32'h5D315B20;
    'h0AF3: mem_data <= 32'h6E755220;
    'h0AF4: mem_data <= 32'h43324920;
    'h0AF5: mem_data <= 32'h73657420;
    'h0AF6: mem_data <= 32'h6E656274;
    'h0AF7: mem_data <= 32'h28206863;
    'h0AF8: mem_data <= 32'h6D726F4E;
    'h0AF9: mem_data <= 32'h4D206C61;
    'h0AFA: mem_data <= 32'h2965646F;
    'h0AFB: mem_data <= 32'h2020200A;
    'h0AFC: mem_data <= 32'h205D325B;
    'h0AFD: mem_data <= 32'h206E7552;
    'h0AFE: mem_data <= 32'h20433249;
    'h0AFF: mem_data <= 32'h74736574;
    'h0B00: mem_data <= 32'h636E6562;
    'h0B01: mem_data <= 32'h46282068;
    'h0B02: mem_data <= 32'h20747361;
    'h0B03: mem_data <= 32'h65646F4D;
    'h0B04: mem_data <= 32'h20200A29;
    'h0B05: mem_data <= 32'h5D725B20;
    'h0B06: mem_data <= 32'h74655220;
    'h0B07: mem_data <= 32'h206E7275;
    'h0B08: mem_data <= 32'h6D206F74;
    'h0B09: mem_data <= 32'h206E6961;
    'h0B0A: mem_data <= 32'h756E656D;
    'h0B0B: mem_data <= 32'h00000A0A;
    'h0B0C: mem_data <= 32'h20200A0A;
    'h0B0D: mem_data <= 32'h5D315B20;
    'h0B0E: mem_data <= 32'h6E755220;
    'h0B0F: mem_data <= 32'h49505320;
    'h0B10: mem_data <= 32'h73657420;
    'h0B11: mem_data <= 32'h6E656274;
    'h0B12: mem_data <= 32'h28206863;
    'h0B13: mem_data <= 32'h203A5242;
    'h0B14: mem_data <= 32'h32353131;
    'h0B15: mem_data <= 32'h0A293030;
    'h0B16: mem_data <= 32'h5B202020;
    'h0B17: mem_data <= 32'h52205D32;
    'h0B18: mem_data <= 32'h53206E75;
    'h0B19: mem_data <= 32'h74204950;
    'h0B1A: mem_data <= 32'h62747365;
    'h0B1B: mem_data <= 32'h68636E65;
    'h0B1C: mem_data <= 32'h52422820;
    'h0B1D: mem_data <= 32'h3332203A;
    'h0B1E: mem_data <= 32'h30303430;
    'h0B1F: mem_data <= 32'h20200A29;
    'h0B20: mem_data <= 32'h5D335B20;
    'h0B21: mem_data <= 32'h6E755220;
    'h0B22: mem_data <= 32'h49505320;
    'h0B23: mem_data <= 32'h73657420;
    'h0B24: mem_data <= 32'h6E656274;
    'h0B25: mem_data <= 32'h28206863;
    'h0B26: mem_data <= 32'h203A5242;
    'h0B27: mem_data <= 32'h38303634;
    'h0B28: mem_data <= 32'h0A293030;
    'h0B29: mem_data <= 32'h5B202020;
    'h0B2A: mem_data <= 32'h52205D34;
    'h0B2B: mem_data <= 32'h53206E75;
    'h0B2C: mem_data <= 32'h74204950;
    'h0B2D: mem_data <= 32'h62747365;
    'h0B2E: mem_data <= 32'h68636E65;
    'h0B2F: mem_data <= 32'h52422820;
    'h0B30: mem_data <= 32'h3239203A;
    'h0B31: mem_data <= 32'h30303631;
    'h0B32: mem_data <= 32'h20200A29;
    'h0B33: mem_data <= 32'h5D725B20;
    'h0B34: mem_data <= 32'h74655220;
    'h0B35: mem_data <= 32'h206E7275;
    'h0B36: mem_data <= 32'h6D206F74;
    'h0B37: mem_data <= 32'h206E6961;
    'h0B38: mem_data <= 32'h756E656D;
    'h0B39: mem_data <= 32'h00000A0A;
    'h0B3A: mem_data <= 32'h656C6553;
    'h0B3B: mem_data <= 32'h42207463;
    'h0B3C: mem_data <= 32'h52647561;
    'h0B3D: mem_data <= 32'h3E657461;
    'h0B3E: mem_data <= 32'h00000020;
    'h0B3F: mem_data <= 32'h746F6F42;
    'h0B40: mem_data <= 32'h00676E69;
    'h0B41: mem_data <= 32'h0000002E;
    'h0B42: mem_data <= 32'h00000A2E;


    default:    mem_data <= 32'hDEADBEEF;

    endcase

// ============================================================================

reg o_ready;

always @(posedge clk or negedge rstn)
    if (!rstn)  o_ready <= 1'd0;
    else        o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

// Output connectins
assign ready    = o_ready;
assign rdata    = mem_data;
assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule
